BZh91AY&SY��(� "_�Py���������`� z�h   �& �4d40	�10��F$�       0`��`ѐ��&��5%<TѐM � 2  s F	�0M`�L$ �hh	��0#MM�C�h�b&�n��D�D����|�#R�E��(¢UR�E�E�'�U~�K�3T��R3T��ғ���
����ЗKW��MY��ſO���
8����hৗ-F�,�E%0��kgk�jd�omR��r�5��s3^��m���nX�9,Y��&םy�'SV�Z���W63ݱfoD'$7�!�֮HrF��&��w�߽˾�4��UU����j}la�>�|�&w��u���J�%�*��K�b�홚��/j�6�Q����Ō�Zٱ���mɞ�Mk�x��Ŵ-�oe��1��^�h�d��p&@��<��FQ%���4�cA�t���r�b��fY��s�l0���m�ў��ɦ��VU*�	�l���Bs�VmVV�Bb�M-�[W���붌�Vlۮ�cL�7˪u��ƒOu]@�!-�  15
�Ҏ����#��>�mS�)JYE�5��]v�ae+�s(�)���TP���u���lD� �RR�CjSm����Y-Ei9ȝ*(@<@�hB�з>�������(d�?/��f�j��,r���^)����F���R�6,Ƀ�Nj��|-v��?+Vg[��a��G�9[]O*y����~�Q�R?8�<���)�Nv��=qN�X|�?��S���~�;$��>���:�0�d,餎(�}kIT��vq���e�&o��$QYe�H�4w��Y(�r���s�x�VN�f��);�RE�2��r��,]��w,�\�ڋ;�>����q��Y���:9R�s�a�=�Nd�Х9$�f�(�\���������(�:$�}���<�����tu�%8�g%���8�]FH�N�c��&�Ga�6t3t��zq�YT�-���E;�W�hѡ�Q���i3u���5:��y�d������Rw)H�f�^d����RG!�w�"��W)QE��9n=�7����ߩ�^��S4ha��Ye���V��r���,w%Ija����-��Y54FK�/��Eu�h��&$�U$��ʜ"7��t�S�p{[���w��9��g�q]e9��֜˺ݭ�}�J��Aa��#EѬ�⊨:��֎S��?s�>��������b9�QKĩ�;T������gS�.��.σsb�ͬ��#���Bf]r�ٷ��389S�ofS%����RYG[��Vni����p]�j���N-o�R>�r9�"��'�^y�j�Q�&�ք�]LN�j��*R8�3�C�N���-$�#cy4�w$S�	B� 