BZh91AY&SY>� �_�Py���������`� �    s F	�0M`�L5Lҟ�zOH     �& �4d40	�11�& �4d40	�11�& �4d40	�10T��Ѣz&I��0�F���Ѧ��I���b�G�?U�`J[��TJ�T��E�'�U�%���G�H�R&VXiI���U*�'w~it�S7�,[��-L0���۽����nѝ+k2S��e�L2�����Juz
�۶�s3N���5]v�r�E�&�2S�pǡM���2�j}2!����]�$8F��M�����c}Ud��UU��Wx�����%P���롉QT斖sd¦~�Ŏ���[Y��.���K���i�������%�3ٺ���|���ܭ)�a�z����e�^�fo+7�U�un��ZlS}2��zt�l0�[/��֍���e�Z֕$�P҂�l8�6�^&EB
&���n����z��)JUpUUUUUURQe���~��<`��G�Sj�s�e���?U����YE����T�жuZ6��4ZҘ���kUI3_EY6�E)�����v���"����:�T��6�^�mp�m}s����o�����i��Y?�����]�m5rv�8���^)���'�F���R�6,Ƀ�N���~�ac��V�7���{�?���<��}��X}��Q��AcЍϝORu7?4��u���Y�7�u�߱E��#�2|�Щ�:ԥ0�d,줎H�|U�MURL���R�>���Ee�m#<�+��U��7.�xY���6�ʏ���-�Wj�T�w��%0ܳ6�af�366����2>F��E"ΖO��(�>���t�ε)�Mfo�FB���0�^�}�C�P���%��^L#�<�������1)Ȼ9,M�e���u�GZw��s�y��������roNT�U%�i?w!N���Z4h{s�Gⴙ��h�5:ݧ��=�J;C7�Iޥ#��m}	c�8j�aICʜL%rR�l��Jq��,dޤM�Qt��u�����jn0�Yb��֏9�m�F�;Ҥ�0�]�h���j���,j�}Mb+�!���&$��S�qN�&��.��}n���}����uE�9�i�u��qNiһ���O9ة#�,<�3r4\�D�ET����`���s�|M&����a�b8#
���S�w))u����r��.��.����F��Dّ��˭3.�jl�����qN���T�V����),�����7L��I�t.��`g�G�7ԩ���J�I�'�/>sTjڲG#&M����jbv���R��1��v򬴓�EIɣ���"�(H� 