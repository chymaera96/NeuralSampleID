BZh91AY&SY���� �߀Py���������`�      �0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`b`�!�24�M#	�Bh�i�G���i7�%w�"�C(��?���$����d��0��T��,�?%���/5H�����2��JO/�+�w�g%��
fͅ�-���S(�Y�w����S�6��ae�)+/C*�U.�wuR�^���u�ݭ��t.�Ce���\��:0��0���64��%6��Ϝ��o�D4k��$:#rx�r��k�˥Y��JU]��w��S�s���Y�V���o�S���]��fբ�=S�li��Ʋ��EQu&ʺ귽[�"6�g�߽��e�O�e��ʙ�c"��0Æ�n��W5]e����KF�Q�M\7f��cʦUU��J�˩f�$қ)��F��\ߋ-�3^�SvN��ֳ߹��ж��Vlf��z���w���U)JR�����������OTx?6��0Yܣ��O���e.���c�ن0��Jگ�^�����UkZ�I�ܳL��ѣ6yk���F1zZ�eH�6�9�l�FKA�CjN��JQ��m���\~�_\�v�s����}Q���],�ϓW����ݵ5sw9%�^)�>�o��ScUJdܳ&�:j����v��W&�=n׹�Ã�}�ɳ��OG�O���D��"��Acҍ�2���o~I���E��Y�7�:]o�Qs�H�#'ĜU?gZ��L��*H�'�ZDnXu3���K,�=�)"��,�FyǕ��U��7��xI���Y���FK�[��X�Ix��RS�3h�va�1ssdY�Q�|�#��A���d�|����a�>�'Jn�R�k3}j2?gy���a���]"�I��K'�^L#�<��L���LJs.�K}�Dsz�:�֞&���#z���ټQ��9ԖU%�i?w1O���h������i3v��$�N�t}~��$����u'���4��K��V�
H�1*t-&��J�7]T�9\{V2pT��J.�]N��{��CM���,P�+Gc9�m�,x%Ija����-��Y54��5yCX���;c�����IO��8�����}N/��}�����uE�;O<��t�'jt��w�)�%I9a�y�Ѣ��ET�h�F#���I�4v86=M���#�U�J��IK�,�Nk�v;��:����۔olț�;�u�e�-M�u5��.I�83d��gK��Ie�>-Y�f������j���NmFo�R~*t:�"���/<��ղ��&N�Iк:ژ�����&T�sLgF���"�U��yT����?���)����