BZh91AY&SY���O m_�Py���������`_z��@ �*   #�0L@0	�h�h`ba"I�! ��    `�1 �&	�!��L����= M2      9�#� �&���0F&
� �222M�@L��h�������57�5�+�H�I$1��~g광0'��>�*0B� ����(��$�!��G����1��:N�<�i�������U���_*I!>�ĥJ�er����mS�f��3ULT�E%a���6��T�(P�h%fPFq�Xł]��tz
�,�鹔�ղ��c[j�6,b;.A��%���K"q����)�n*��QQ3L�"�F���63��TH�z�H:���$��ӹ����t�(_�|`� Kl�،ہb���a$�35E�QcE��!�/�x��>��(ެ�H��Z$�F,�G�_BM%�r�#X$�'��H�ia�s���d�!�td1�:%DP1� �]�q�A�g�� V�:���:qH\4�(6l� ��I<#�R	�d�e)��\SgF�%��6s��V��&0b����TI�ƫ��3D �pBۓ�����ppIl�c�h��j�5*�@�vL,�@�A�V�o� {��v4�*x�V͛-��:n�!V�Y-�bpQ�4QEj	/�ǥƮ)̹���Mg��Y��2����Ll�pL���GBb�`l`�\IF}+�"՗B6���lUUUH`�$���������x*jS�z,��Qg갘.�S,�ʱߚ�֡1�0hc��@YC S���$D)h���ʈrD�L�����cHc7F�һK�ġ�����G��T��od����q<_�q�����"����0|������Ӫ�܋�����[���&�B�1iY��Nz����v��F�[�����ڒ>q����O7Ğ�<�H�<j��Z�kyT��C[�L�)�R��$S����\�${bF/mT�8)J`�b,餍�w���UU!Q��=��YgՓ�0RE�93������TY�u���:�楘�ԣ�,XY"���NJ1RE�(2���fL�.�fř�Z�gaG{�1<"F�5г���pܔtc��I9�O)�&���s��0z^�|�[\�I#7	,�r�`������8qL%7�e%���b7�}Fh���K�ޞF���#�i���7�&��E�Ib��ݼS��~vlٞ�z��-&N&�2S��H�zd�����ܤ�R���5<�cs(hi0RG1�;S�i$`��JTQ�ꢛ�=��*@�%N�΂�}B�#3�Y��,���V�����R2d��D҆QB��dP�FhV-q#���\w�1#�z�$�
�S�nM�M��]'��m{����v�:"�N�u��nN)λ���O9ҩ#�Xv��њ�#D�䊨8���H�a0?�nN�7ScQ�k��a��TR�*uε%.����,�r���/�[J�mLI��	�u�SN�������6��F+-g;kiIeX-���35I#��w��s�M��6Oj�6�)��T��G�Yy�0:#CR��F,[��#�tph0��k�Xґ�0ʌϥ:Jv���Ƣ��-�����"�(HK�q��