BZh91AY&SY�� �߀Py���������` Һ    � �`�2��j�jML�C#h�4ѓ@ ��0L@0	�h�h`ba��(02`Li���	��`�1 �&	�!��L����M44di�4�����M�݉�-)�?��-R�'�Q�D��$/(�������Iy$�R#�H�H�Ya�'��\o��ݤ]-^O%5f����kS(Ⳳ��Υc9^�م0QIM��
s)��T�?���u���צ��6���l7,e�Y��6=K�p�MZ_*5e�5�^�9!����W$9#bx�Uϳ���ۺ�4�R�UWk�]�:��Q��S���q��K'Y��)�aJ�Ngfȶj{Xi�c>�6�U�Z�|�zmV�mae���m��<��.B����d׊���S�����l������㙖|�0���,���ٺ�e����UY�`�YY2�Gnl�H�%l�J4��͓
�������/�ꦁBI@  a�����j��;}ڧ��)e~�G�u�Xa��X��F�F��f�MYL�X�����=�p�=�d3!
0���ػs%�ȡ�'#�N��R�ԛv�w�J�)�|����(�pTQ�r�	��q�X�K���S��/��UJdس&�9�������Xz]oK݆������=y>�t=��~Qh,z���S�Nv��=�N�X|�?��NgC��\�>���N
���JS�BΚH�'�b�R�
�vq���e�6o��$QYe�H�9��r�d��ˬ^�s�y[VN�g,v�S%$]�!IL7,͢��Y�r��͍������I��t,�d��G9�0ޞ�'2l�R��k3|d.~��[�����*4tId�����O|~��֘��]��&번����:�Н�&���F�Ga�6t3t�-�Ƣʤ�m'��)�ڿ3F�r�����7Y�R&jt;'��{��t��o:��JGK4��%�Vpհ9C�9�%qR�Y�JS��ܱ�z�7IEӿS��'Ȧh��Sq�0����h�g!����Ѣ�rT��K��к�U�SI�Ư�k]|G\���$��S��N	7��t�C�p{ۇ�l;���t���8����T�Ne�n��='J��Ya��#E�'�*��{�\�10'�r�������7G@n�DaTR�*v��%.���8�Y�싨�˳��أsk"l��deЙ�\�6m�k389S�of�VKS����������CEG��w���q8�xپ�Hp�)��T���<���`�[VH�2d���9GCS�ڰ�ɕ)Sѡ�IN���x�T����?���)�`