BZh91AY&SY2+� �߀Py���������`� �    9�#� �&���0F&9�#� �&���0F&���ޤC�       � �`�2��� �`�2��*HA��CS&=A�����SM�݄��Ȍ�H���`����d��0��T�Eҋ*O�z���K��R#�H�Q&VXiI����[�v�h.�����ae�~�5��qY�w����Ly4��*aLRV���.�L���S��W�f���ft챼ѵҺ�匣}�5]��l�pu5���k]*63ݢ�<���hHfƕrC�5Oj�����6�f��(UUv�U��O���"�*�W�_U,�f\��TǢr�'ģ��g��T]RZ�|�����m�����^��y[{Ɨl�X��f�6�VZ�Y�w��ƌ�i-fkg�~E��3t��!@(:���[i�h�D"�c�4���
��e5�w/����s��ե�7Sf�T�����SÅ�I�w*��)U�UUUUUUIIe��;��c�v(���S�)J�Qg괞u�ma�Qi_M�����K�V��/�YJ�*��{ڮ��j�j&�X���Jm��ڻ6KA�CZNG�Nz�R�n�۵{�������k���g#�m���d�|�_���f�j��,r���^)�~_M��UJdس&�9�������X{]o[Ն�	>1���y��'��j<*O�-�27>�=)�����)Ћ�g�ܔ�t;��E��#�L�RpT��
R�E2t�GY>��Mb)9�ǻ�K,��{RE�Y���N���%n]b��NvOj��Ŋg-ֽ�
�)"��Ja�f�.��;�f.lmE��G�d}Sq��Y���:9R�s�a�=�Nd�Х9$�f���\���w�����(h�������Ol���LJq.�Ku�Dqzz�:�Н�&���<M�n���l�f�N-�ƅ�Ib�O��S��~f��}Q�-&n���L��v'��z�t�Fo"��JGK4��Vpհ9C�9J�*(�b��-ǭc)�R&�(�w�s�����jn0�Yb��V��r���,w%Ija����-��Y54L�5x_sX���:������IO�8A�}ˤ�����|�{޳�.��y'�S�ʝi̻��ا�t�H��#r4]5�<QU[�:Ӕ�`�߹ʟCGS{i�n���1�¨��T흪J]aejq\���QїgŹ�F��Dّ��ˡ3.�jl���389S�o�����pp),������74��C����s8�Z<,�r�8}T�s�E�>�y�9�VՒ8�L��ZE�����v�>�2�#�c:4>T�)޲�O
��67�G�rE8P�2+�