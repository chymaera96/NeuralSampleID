BZh91AY&SY��M �_�Py���������`_"��    ��b�LFCC �#	M4� h      ��b�LFCC �#O�H  �     0`��`ѐ��&��RI��ddd�'�`�d���4=F�F��oRl�I]�I-$F19���K�Kx,��E���$�"�*O�~k�U��	��G�����a�'_ګ~/'vrF	�]��F���o��.���-ʾ�m�3��1b�uG$!��^4V%%2�x�6��*#��L��.!�f�P�\7�,A���@��F�
f}��
�j(�i%��
9%I4�; ��\f�S-w$9��&�w��kU+�"�*���q�O.��}���	Ļ��k�����Y��^�[�_&Ǚ�l���! �  N�13`F]+eN�d������J�}k�t�cJ%1��=V�؇M����0�!�A�m�u%�ѩ�z���J��"�Bxx�-�w�U��q0Q���H��ܚZD�w�p��i�|t�-��Q�˚�OKaP�=0E�zҬ�x{Fq0ȓ7�I0"8*vⴱ�NFK���Z�5�UC�vI��������@�!!�  0bbi4�,LM�6��.Y�G�����,���i#���Z뮲��0���dQiq̔.�.*C��2L��C�:L��j�Jk�b��4b�(gI��� �I����ym�x���Þ���1&i����������]4or,nL���}���D�h�LZ�b�اEU}>V���ӹ��{�����ڑ��n��=x�}���r�?(�=(��)�N���>ȧX}?�Ȋt8;_�F)#���M�������LE�T��OcS�*:YG�饖}=˩"����YDw��T�TY����'K�ֲu��(�NEJ1T&$�J]�fL�0]eݫ2��giG��1<b6�BΆ/!�rQ�}e���t&�
S�M&O��F��.�=��}��B���$�z$�<㽋��p◔�`�Kfb7��e���;K�O�zy[��!��'TF�2o�"ʤ�l���)��á�6g�G��-&N&�)��#��=�J:�S'�Iڥ#��k}ics(h�]I��ޜ�IJޥ*(�R����c2�F�(�;�:L ��e2Fe��u�X�?����C)��5�ԩ-K��=l���F�š�F+;�kH��q����~
�S�nM��a��O�m{���w�:c�'�o`����:8���J�=E�{�،�Di"yb�/h���EϽ�������k=m��6�:.�)�J���ILV���nQ����65(��Ě�911��0-MZ�ZDdmnM��ȥbt6���Q�sɵ�'D��RG����сq�M��̟j�6����T��?��L'���5���#.f�rG;ph^rv,<1cJF��Tf|��S�e���*H��&o�.�p�!�