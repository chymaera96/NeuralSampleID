BZh91AY&SY�zD� �_�Py���������`� �p    ��b�LFCC �#Jm1�@ � h    5)���<Ԁ  �   �O�T�@  �@  � 0`��`ѐ��&��RBd��	��aM4��z�F��m&�I+�	h����G�?U�����d��0��T�E�ʓ�^�����"=�Ԓee���?
�W��ݜ.����3xYbߧ�ja�Vv]����)���f��.QIW�g�)�S���N�9]���\�fi�c������nXȫ�h��%:��y�s3b�n���6.�$p��C{\������=��~�ͪ�5��*��_��֧�F�FJ�f��m~U%J2�Yw]VY4Vk3Tc��ֺ_Gf��ֿm7#}DaKQ��|�Y�o��ZpT��7i{�[Sa�3emo����pa��U�-h��#m�l�lݫf4[�y�n*��u� (����(N�a 5��,T8j�d�-gQ4��A!�XTQ(��`Sf��I �	Pi!��/!Rb*$��\TP!B�   R����'s�ny���>�mS�R���?U��.�k0��++�4`��5��1Q�KT�mj�Z�e���//JU+FWҖ�ک��3����2Z�i8?�x**��u&ݫ��o���?ݮ�v����m?�C'��j��>��m��.��:]�������Ѫm5T�M�2`�S���]����Շ���=os�s���"y}l>�ya��*O�-�:7>�=I�������g��%:��آ�d��I��NeO��JS�BΪH�'ѱ�/H�T�,��祖|ٽ�)"��,�Fy��s�Y(�r���:Y<M�'yFŋY�Z;��.������f�b�,ùfb���Y�Q�xfG�MŠ�Vt2w�\�GI�0ޞ�'Bl�8I���Q���;L=l?/˙�(T4r���/&�6Ol��֘��]��&번��w�98G$�16?�-�;���7T�[ӍBʤ�m'��)�ڿCF�Z���|V�7Y�RI����{��IGS�f�);��u3M�*X�g[)#��xӂ��W)QE��9�=k7�$�%O�Ix>O�Lѡ���
ae�)�h�3��F��h�c�*KS%ޖ�h]F�ɩ��,j�>���u���&$�U$��Μ�o_r�>�������x���1t���8���t�N��n��<�R��Aa�y���k"xb���u��bL{�9��h�7������#�0�)x�;gj��XYZ�W,�;"�9e��nlQ���6dv22䙗\�6m�k&g3�9�{5d��gC��RYG[��7D��P�9�{ڮ`g�G���T�7�N�H�	�Kϰ������L�7����ɩ���X}2eJG�th|��SƲ�O��67�G�rE8P��zD�