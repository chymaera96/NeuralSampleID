BZh91AY&SY� � f߀Py���������`���(�   `�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L���HM4��ڀ�  4 � �`�2��*H� L��CS4b�=CG���3SM�لEwI�I1���G贑����d��0TJ�PKĢʓ�^������"=T��C,3����[�o����$�][##qA�/�h�A��	>�,��k8�F
X���m��ާN�Jq��ܳ�w2����ll`��M���\�އ�_~k)Q:ٙ��6oQ&�m�H�SV�$7F��&��w�۵�b�M"R�$���M��� ̡9�$� �2��i&Ԕ#X:�U�G��F��B¥����t�饢��cn��g.�$1Rd���R^��A��o�R��U���6�7^�a��e�8q�D�e&cTo��4$$XȐ�L�U́�lOji:R��0���K(&�%E2yo��P�YP�R�3��djJ5�<fd!�j���*��dF�&�j���
2��X��h��y�u6�q�"B�%�I$�I$B���9K��(�DaOAJR�,��z�]��(�Q��s;�I�����b����[v,I%�UA�DFV8��0TpA�F��� ��"1�d�-�W7��|��|[������������Eڵ�G'B��k;�=����͢k4T�-K1`w)ƪ�?���X��у�v�of��>1����'��O���<�A�TO�-�J6>�>��l~I��E9���,��"S�����\�$}�1}	�S�sR���Y�I�d���Լ:�G��K,�پ�
H���&q�Q<�X��b���u1yZ�N�2�b�Съ�x��RSř3X��;�d.jkE��7�b}"l-j�����(�<���qM\Ԧ�4�=�1?Wq������7��$��K'���#�<���S�ja)Ȼ),M�c���9�G4�0��$�6-�:#W6N���S�I,�K�~�B��k�f͙�Q���i2v�*!���"{�'�IG[�d�);Ԥu�Mo:X��5)#q�<r�L�)J�,ԥ)��ر�j�$����^��S$f`��`�,�A�֎�RH�Fl�;Ҥ�0`�z٥�u+�q1X��}�"+����=fUI)�pM�m_b�>����lQ���ꋤv�i�u������wk��OA֩#�Xx<͈�x�H�H�����8D��߱�>fn�ֳ���`�7#QKĩ�;�������gc�]G<z|[�lkbMX���L��Z���4����7��LV���-��%�v�<[�2q���I�o]�h���'&o'ک�E7:�"���}R��0:�F��9Dŋk[9&��͡���X~���#�a��*u��Yi'�EI�I����"�(HN�� 