BZh91AY&SY]��� �_�Py���������`�      �& �4d40	�11�& �4d40	�11�& �4d40	�11�& �4d40	�11�& �4d40	�10T��L�Q�d=L��zji�&�9$�|Ȍ䆲?C�X1	K|�O��
�UJD](���W���$��">�>T�*$��i=5�V�W�At�YgMfX�ˊ��
9�����z��^���0��)+��ώԺ�Ju�
�Y��s9����#{s��oX����4V64X�3-�^F��\�j���p�{�"C{n��$8F��M��o���UV4�
���~�<�j�5��q�����e-'2ו�`�h�S/l���g��)�T�"aI�K+'ŕ�S��T�W�+���}I���7��f�l�س���6&i����fشb�^�]��b��^��*p2m��}�Cѽ�U��V�%�^���kd�ZU_~���_�9���۶g�ۥ���.����<UJR��ܪ��������*{S����gr���j���e�]E���]��0���<|�[)���
͵���ĵIU++Z�_,[���ک��1=ͫ�2Z��p$�R�R�ԛv�v_m��6�g�5Ϟ�wS��8S��2�����l�M\�ŎIv���}������6��S&ř0w��U_/��l,u�j���z��7����&�cҞ�ȟK����?X�=���)�N���=�N�,>E��)���~�;���2}	�S�tR��)���I�Y>jة��R���}��Ygɛ�aIVYf�3�<�'*��Y�u���g['�ڳ"��j�l,Y�T�RE�`RS�4h�va��\�ڋ<J>o4��&�Eг�d�:rJ���a�>�'Rl�8I���(�\���[����.�B���Y=e��=#���G�N���Ne��bn�(�owa�G�&&���f�Gq�l���M�Ԝ�YT�-���<[W�hѡ�Q����f�9RI����{���#�f��<T�y���K��V�
H�bt��W5)QF˪��+���M�$�%O>�Yx>/�Lѡ��S,�P�գ���d��,x�Ija����-��Y54L�5y_cX���;S�����*IO��8��}ˤ�{��n����qt���9���NIڝK�]�z�"�����-��t�D�ET���NF��I�4v7������#�0��^%N�ޤ��V�5�;�uw~m͊76�&̎�F]2�ũ�o[T���S{5S+U�gS��RYGk���Sө���W~W03�ͣ���*C��N�H����/=�յd�i�&�փ������w�>y2�#�c:4>4�󬴓ʢ��������H�
�]~ 