BZh91AY&SY&#[� ߀Py���������`� w��    `�1 �&	�!��L�����Q� 4  4  �x�S�4        Je$�2h24�4�i���h1� �`�2��*H� ���2OS L)�A��Q�=4M�ـWb�1���~�!����d��0TJ�T���ʓ�^��Y%�d��d�$���;����[���f��mwcM0Yb���0`��λ�_��ٳA�51R���%�t�L��S��Wb�|�e26k���[E�m6,b_u�)��L�YO3J�)Yx��ˬ�����I�rՁ!�.��s��4�)X&B�*����㚟E�E7׫���eә��U�JV��D�uj,�+,��h�U�6)r궧�i6��R�?��^lU�h�Zԧj�����Z��u���N�!B�NI�d1"�LC�����$�!(qBtŔ�Z-2C�m�Р�U$�aqVH�^��
f����VJE���0�}X�ojn���%m͵���_�&]���UJR�%�$�I$�! ��pMR�7J>�kS�R���?E��]v�,�`�I�$�����5�)�MI��!�ԭ�d�Z5�E)��g��vLV���M���)F�Mz׻�[��_L�v�����n{����/�������ծ�8�����?/�mY��1jY��N����-v��O��7��������x����a��ȍr���Ǚj���l~i��rE�̳�l�rv�b��rG�1}I�S�rR���Yऎ(�}��E�K(�y�e�6Oc$QX�8�!��p��E�X�?��b��N�2-�T�lVH��"��6,ɚ��,�ڳ!sSZ,�(�<S�6�5Y���9pJ:O!�j{d�	����&�'�F"���0y��~_��@�H��K'���#�;ؽ���.i��줱6]�G���ɺ9'i���S�ض��<&�L�ŵ8�,�K�~�"��k�3f���������@�NN����%���Rv�H�2Mo"X��5)#q�;�r��+�����JR�.=k��$�%N���|�"�#3��0Ye���-L�2��0�٬v�Ij`�.�3KB�4V-�+;�sH���s���O�%>��!�}��������~���Y�H�x��S��9�B�nƥ<��RG���x���I�Psz�1��`}����C7SkY�l�A�a�����T읊J]aehq\���Q���cR��lI����$Ⱥ婫_KA���7��J�V�t7���Q́��ѓ�ff�x��{�.`2�ś���T�����*�H�헟i��5���bŵ��7.�M'[�a�ō)S���S�S�e���*H��L��]��B@��od