BZh91AY&SY��K� �_�Py���������`� �t    � �`�2��j�j4�=FM4����`CA�@9�#� �&���0F&���        `�1 �&	�!��L����L�`�54�4h�4���3D�M�I]�,��!���~k��+'�Q�D��B.�YR~+�W�$��"=t��ee���>*�����]<+����Yb���Z�aGR�����cӢYl[
`�������fjf�}R����4�\�fp��ѹ�u����j�f�ۭ��_t٪�Ū���)�,�]��v���/�	h�;�Uϯ�o�p�Y��JU]��w�ا�F�"�������,��K0���{��^�9�{˷{Z�-��v7�U�Z�O���p�)(F�3�>�~���5�{\o�*����Yi8Զ���ͲZʽ�gim*�Usm�-z�4��J���ͫE+'6�LTΛR-��L��&�V+
�Kf����>��g	u�Mr�3��^�-&�!BH   LM2�ck�x��;T|�ܧ��)e~kZ�0�(�Y^�_M�%T��j�Z�PeTUjVՓ5�eR�7*E)��O���얃"�Ԝ����U)F�Mۗ��"p"S%���̨Lj@P �QDCXM��(�r�ic�]���c���:5Mƪ�ɲ̘;�窯��k�,trj���z��88��Mη�>��+�8�x)?�=H���������)ԋȳ�oJs��W�Qs�H��'ȜU?WR��L��JH�E���#e���>�U,��h��RE�Y���O�VJ,޺����C'��d�Q�ibӴ�j�RE��d))����X�0��\ٹyJ>/4��&��h�9�;ήIGA�pOt��6�R��k3}�2?Wq������s�4uId����Ot~��ؘ��.�K}�Dt����4u'�����S�޶��;ͺ������4,�K�~ΑO+r��4=�;:��-&nÕ$����O��{d�yc7�I�R��f��:X���0��c�Ne��T�El�)��ڱ���7�E��S����h��Sy�0���u���F��h�cʕ%���cD�.�Ud��2X�����WgH�O��1'�T��w$�����}�/sx�͏ڳ�.��z'J�)�䝉λ���OI�T��,<^��h�k"y��Ǵv'#	��~�$��:��c|u��FE/�t�RR�+S�rηl]GV]����7�2&�����2떦ۺ�g$��%��9�\JK(�`��՛�hh��q]��\��'KG�7ԩ?%9�
�C�O�^|��չd��ɓ�sA̺:������*R:Sѡ𧐧��I<T���4�w$S�	/$��