BZh91AY&SY(�0 _�Py���������` �@$*    � �`�2��� �`�2��� �`�2��Jd)��G�4� 24 2 P�0L@0	�h�h`b`�$�Bb2=ъhѣ&'���Sz�e�Wa�I������^��,��E���L!(���XUW�$�"d���I��ee���o'���ߣ�ݜ��yk����.�ž;֥�Q�gf��+�#m��t�KRR%�e1S���NI]�3ご����f��`��sUX��V,�����ږ�a:Y����Jz�m�:`DMM/�rClh�������t0�db�I%�<!�� �D�Z;<}����,%nm��URm�,� fx)�#LxN��0*�[G��ҹ߉������g�����EQu%�����bQq&9�)u1�'�g�L�4�3�!((Z\��t3�;}}J�������1ˋBޜ筁(�0�+��,���K��E�cu�U(���:�,Wa�E��Ҋ�4�+yf��A�A��y���I!VEƧosh��a��jp�\Uc6�D���.v�N��̝)��ppt�-�b原�c�=�#��!/9UUUUUUIP�eO\'s��xE�9(�S\��JT��?e��0`ֺ묡�����4��Dn%@��7�̧��WE�Qd���X�0Q"BH@�(�E��F�!Aq�6I�� X 4��>R;�	Dr��ɒ����r���ۿ������b���??�ŃV�h��Xޘ9���nӿH�dP�42��zK������.�u���w3r'���O:z>�x�}��H�"�?X�=(��)��Cc�K�TS���g��	Nws�Q��H��1x�r���JR�"ΚH�"��SSKQ'C(�zie�O�u$QX�8�(N��}V*,��c}��kY:��L�,ZYȱjIɊЗv�����d�c�]ܴ�`jkE��'�bx�l-j��b�8�J���]̞�':j�6ɤ��Q�����Ol?��(T����O	.�8�b���z��Ibl��G��]Ŷ8�qy��8'��m���5qd���I¤K*�ų�À�s[vlٞ�}Q�֓'Y���)����=�J:^S'�Iܥ#��k�����4j.����ޛV�.��JTQf�)M�b�3�I#d�`��|�#2횊.��Yb�?����D��٬w%Ij]t��f��
4V-�1X��}m"+�������}�S�oM�f$�=��k`��G{޳�0H�<���oN��`�v5)�t�H��;b3a	��动:���	��%ϵ���f�s5�����j.��a�d�RS�����gS�`��_�cR��lI��)���5k�i	���7'4ɍ���s�7E%�u�v�f��<�*D�s���(����Z�7x��Щ")�O1s�4kY#�&,\�l�M�šy�ذ�bƔ�	|���S��z�I<�*H��&o�.�p� 8Q�`