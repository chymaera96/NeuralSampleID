BZh91AY&SY3�Z� 5_�Py���������`�zP�
 P   � �`�2��� �`�2��� �`�2��I��AG��2�C@  ��0L@0	�h�h`b`�"�224L���jh�i�m'��M6�n�-	1�����h���+���*$��(d�KW��\�d��d��a�'�g:ޫ{�O�];��hт��������+;n�{�]M�u��'��0$m��\с,N����ܳ��L����Y�5�n6�b_���
S�-����(�W��u�0_+.��D膶X��D]<�������סY&�)B������9��Q��)�Z��z8ү��hOP2�ɛ�ș(s�;�ǸՃ�Mu3�־5)�n�T`��K�U~�x��K��)u֦�c�L`�ҷ�1g!�	�!��֋`�z\���M������J�f�:ި�#�F:��YYк�4Ҩ�e�2�R��a,0`ڃ��ro:g\n{Vl�н/;nkfe��V�b������N��>E��3m{k�<�׿���w��UUR2T��w����a���C��=)K(��Z'�uڰ`�e*ؾmJ���)A#�8�����KUK-$ة��'i<F� �7I��d�䓎��������i�~��C����b�|=�g�v�i�����.���O��q|sh��*SŘ�;�骯��k�:�4`�9�N���G�Ǚ<�y>Vt<�4
��Š��F�ΧҝM��0>��$X~���l�t�;߱E��#둋�Mꟳ����"κH�'�w������%~�O�$t�&q�R<[�X��j����L_3U��F�X�v��Q��.�A����2f�v0w��\��w�|^Y���t,�b��%G���=�N���JtI���Q���;�����{�P���Id��y���?�r�Jq.�Km��q}=�N���c�qO+j�c��92u��ܜj%�Ib����S���,ٳ=j9�Gⴙ9�*A����=���$���2y���R:�&�:X��6)#��)дL��J�,إ)��ֱ�r�m�����Qx>�L���Ci��,��$�+Gc)�kFl�;Ҥ�0`�}�к��C9�h�}m"+��G��$��S�pM��ںO�������6/jΨ�G3�8���.	�:Wsw6)�:�$z����#I�Psz�9$`}����7csS�m�A�a�TR�*wN�%.���8�Y�틨�o���F֬I����$Ⱥ婳^��27�&���Jb�t����Q́��ѓ�ff��f��֋��qf�d��!��C�R*'�<����Ѫ�dbŹ�8���C	��X|qcJG�*3>�)��O$ln&o�.�p� g�P