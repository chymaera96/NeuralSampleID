BZh91AY&SY��� �߀Py���������` O@    9�#� �&���0F&��FP �     `�1 �&	�!��L����   h     �0L@0	�h�h`b`�!� MM14"=LOQ�L��j8e$W�$��9$k#���p�	K��?Ҍ����Ē�T��U�d��*D{i)!��kI���+�W�1��'�z=��d���?E�&J9����Յ=z#
YE%E-N*x��)��+̶|�i45�����B�Λ�l�s��_Os�sY'kq������0�ȑ�z�Ht���MX=��Ã^
�6�R�UW��a�;����ɾ���������s�L���f��5�Z�k����kmY5Tk�i�Y���f3ݶ��	�Q�3݇eRI��Ij��Z�����o�/����O�Tt��i���O&ReT�V�FVt)��f�2��N���2��)��XՕ�Z]HA��'��6�ӄ����F4�b�H
�M�J阫1�����Vf�1V�7��2��ݹ�m�SeU�i�����u8W
��i;��-)��!$   &cM2̓��޸ȷ��������-E�U��a��L�-E���Q�.�kwUwuR1Q_�£:�6V�F���[I*�z�R���}M�5f�3(n��	�U)G
M����]?�񶟻myo���/�2o���������a�}6rxqL:�)�?�'�Vɼ�R��-�#�N���?�qgg̞�{����u�[��R}�>V?�>�6uI?8�,�#��S�N���4X��	%:��Oأ���I3|�ԩ�9�Jd�f-�I�i�k{�;G�쥭�5{�)"��=ƚI=.��Vj-������3zӹFM$�\x࡚��<�f))���5Y�Kd�[A�sz-�Q�z&g�I��5U�ټ�>)Ga�:�u��jS�M���Fc��2{_l?���u��rZz�I�=C�����N}锧#$�p�8�O��������n~I�p_�<��m�NN��PZ�,�g��)���[V�O�Gt~+�GyƤ��sxI>�a��(�z�'���։��%�ZCf�%$t�Cҝ+�$�JR��nR�����Ш�	(�zv;A�|
h�L���kYHe�sI$o��V�<���d�0�Z��
6Vm�d����}��+���{�I���RJ|�)ԉ��|����\�n=/�n��GyꜘZ�n)ޝl;�-�z��I�ǥ�pF�I6�=U{��N&RL����)�5w:ϥ�9��t�%QLD��<T��ūc�������\�pofMٞ����.���6�hu8�Rt4f��n�S����7SV������:�}�2D���h�!��S�ة�O�b|�Gdl޴�RLٺ����9�2���6t�rL��S�NҞ��I�QRF�A5�w$S�	�y��