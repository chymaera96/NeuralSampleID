BZh91AY&SY%Ul� �_�Py���������`� {    �& �4d40	�11�& �4d40	�10�j<�� h�     S�T�        ��b�LFCC �#I#Q��z&��LF���Ѧ��I�"W|�-$2�i#����L	K|O��
�UJx�ʓ�^����3T��R3Q&VXiI���\o����K�+Jh�0�ſOz��
9,���h����Ш(���t�=
w��)��+Ƴ���s3m�t��]�б��;�Ռf��c*zXY�;Y8�FoQ0��ѝmrC�0�4�s���lߪ�Mb�*��ߪ�!�O���"�kz��YIۗ;K��\Ɋ�h�S?\�f{YM"K)7)e{����o��v:'Eow��WȘl�Ukd�n:[i�u�wj��[�h��k�{,��UoVmغ�]����Z�{��:�����0���
hk��
0D6�h#E,2EH����M����$�Jr!A   	�Zz���4|т��M�|Ǧ�)u~�&]��0���᝴l���)v7�^�yj�ij��VW�U�j�z��*7�E)��Ocz�-Ei:_�9�)Fԛ��w�]?m���]9o�u:_\a��멓��j������髓���.�ix���<���UJdܳ&�:����Z�Ŏ�-Xz��׳��#�{���'��퇢MG�Q�Š��FϕObu�~i���E����m�v<�E��#茟pT���R�E2v�G$Y>�5UHRu����K,��},)"��,�FyǙ��U��6]b������oY�%.X�qFJH��B��l�6�af377�����2>1���Y���;8�g�á>�'Rn�R�2k3}�2?gy���C���:�
�Gd�O���G�y�>�����1)Ȼ9,M��#���0�t�bx��s�y[-�w3wc7lrt'*�ʤ�m'��)�޿SF��G?~I��ƢL��wG��>y%�)�Τ�R���7�	c�8j�aI&!�N���W%)QF몔���c'B�M������/��)�40��Ye�z��g!���ѢǂT��K�mк�U�SH�cW��5��|�8��f$��S�qNоˤ��[��l>�q�}�:���<��u8�4�]��ܧ�v�H�g��4^5�<�U7�9���~��<N����;a��FE/�|�RR�+S��'t]Gf]߃f�7�&��F]��u�Sv������8'C5R�Z�N%�s`��j��44T�w�cU��rh�3}
���S�֩'�,��Lq�z��&N���t��Ʀ's�a�ɕ)�ѡ�iO2�I<�*H��&��.�p� J��$