BZh91AY&SY���� �߀Py���������`zqͶ�   `�1 �&	�!��L�����DO0��@0��9�#� �&���0F&j��z�4       � �`�2��*HB��#S4i��A������4�M��+�I%���"i#�?U��R�*��!X�* IHA
�OB���)f��f�FVXiI���ޫ~.�6�E�*��M�,�o��0+;.��:7��v��t�asC�dY��tM�-hO��"�;��uw�vG6���vp�66,A�a���0��ɓ���Q/�޴�a��ůz�h�L�F���47Y ���w$9�ZyR���7pnެ�TE(UUv�U��Z�*5��s��q���	�9�勊ɤ��]%�~�V�صz����!�'�.+<o}#��9�r�r��JJ�4��==���FZ�)�p`����ͅ
�`�>7T0	�r��B�;W<C1k�Au�>Q5��!6[E�Q�zx��X����Ú˳F�Ǵ@c,�z� rV��C��1��r�>{n�O��I�E��t�򴖪n\wkE%b�Sr���h�g�9��|2؝mg"ռ�[�*w	��ы�=�,��:���g�"".(�����,��Dw?FǦ0Yأ��=%)K(��Z=k���,�ҭ<t[j��D&ID��C��☄��209+A�6��B���R�.�%�-K틴d�6Rs?��ʔ�m&͋��~���yX����p}�X�==���(�x���qv8%ۚ^)��/�a�R�5�Ƀ�Nz��|-v��G��[�z��ޑ�����=y>vt=F�ި��-�R6��>��m~i��rE�ȳ�m��;���\�>���2oT����0�d,餎(�x��/R:��꥖|����Ee�m#<�<�Y(�j�����fœ�F�-]�E��ة��0�A���Vf�b�,ùfb��Y�Q��̏�F��h�9�<�.	GA�0ܞ�':k�9��3{�d.~��[���os�$h�%��^L#�<=��S�ZbS�vrX�n�#���0��I�bk}�)�m[lvC_&n��-�Ƥ�*�Ŵ����sb��4=�:��ങ��3S��#��=�J:^S7�Iܥ#��lz�p��aI�!���IJ�*(�Z���j�Mʑd����/��)�40�m0�Yb��+GS9�l�F�;���0�]�h���jVMF�,jw������:�>��ğ�RJy�x7/�t�3�o{�G�k<��t���8����	֜�ݭjzN�I����mF��j�<�U[�:�8���?s�x�:��clr�̌*�^%N�ڤ��V���NȺ�Yv|Z�mldMy���&e�-M{:�37�&����e��oo),���ɽ���hh�#�޻�Թ��N-��Z�7���t*EI�}��0tF�Œ8�dɹ���̺95��Շ�L�H�΍�:Jx,���EIۉ����"�(Hv�\׀