BZh91AY&SY7abq �߀Py���������` ��   �0L@0	�h�h`ba���=OS 4�� 4�   � �`�2��jmJ=OS@�       9�#� �&���0F&
�A M�jh��'�OT�i7`�ڒ,C"H���d���Y?�*%U*H\�ʓ��Ū��5H�U#5H�Ya�'~��+�v�f�K����6X���Z�aG:Ϋ�_��:�]��y��K�RVYgn\2S
vvR���+�f�ng36kcyu��]��c#~w,�&���OK&t�¦�m�0�HrCm�!�l�!���6.}��]�]�Y��(UUv�U�3�O�Mk�q�*N���xf¦������l���`d��E�|�]E+e6��.�x��k>��i�lef[A�HN$GJ���h�����K�E4�=�Y��/)���7�n�eM�ے�^��m]�9��~r��:״��r�JR�[ꪪ�UUT�Yi�;��c�,�b�}ڧ��4�"��,a�����ma��.��r�4�̞�dUg4ƫR�1�d�k^�dSZ6�E)��cb팖��'�h2d�a���鯞2'�L�*�<.2���9�?�3W��}l�M\��d�{K�>����Ѫm5T�M�2`�S���]����Շ����xor��9�]O2z>�},>�y�Q�Q�Š��F�Obt7?4��qE�̳�n)���~�;$����'*���)�S!gM$pE���إ�R�Q��>�M,����0��+,�i�w�y���Y�u���ΆO��d�u�dбn¦JH��%0ܳF�af�366����d}Ť�*Y���8�%��z{�鳊��Y��!s�v�z��|W8�I���OAy0�0�d���N=i�N��bn�(�gQ�$qN�c�pO#rۣ��8�t�Ӆ%�Ib�O��S��~v��}Q�-&n���3S���zOt������Rw)H�f�^t����RG!�w�"Ʉ�
UUY�JS��ܱ�z�7IEӿS��'Ȧh��Sq�0��'�Z:��g#lb4h�ܕ%���[D�.�Ud���cW���������f$��S�s',�z��I�>�+��>�a��,苤u�i�u��s'Zs��v�)�:U$z����.k"y"���u��s�9������zۣ�n�DaTR�*v��%.���8.Y�싨�gŹ�F��Dّ��ˊf]r�ٷ�����NT��YU��s�\�%�u�x�Z�s��g*�U��ph�}j���)��T�O�<���`�[VH�dɽ��r.�-LN�j��&T�pLgF�ʝ%;�ZI�QRF��h���H�
�,N 