BZh91AY&SY�=y +_�Py���������`� ^��   ��b�LFCC �#S	����   h    s F	�0M`�L5?UC@ @     �& �4d40	�10T��h���L�F����h�I�Wy�$F�?��,F��'�Q�D��D���*O�I�1UWHf��f���JO�%qU���B]<Ֆt��ae�~_���
:Vw]��4mS���F�E%/�����\i��S��S��W�ξ˙���69ۘ]wz�G.7,ьlh�rhYm3^��jj��&�OT'gh�oc]�$8F��&�ϧ�����Y���
�����v��Q��S����I����������.±�Yo\��B��^Ƙ�Y���R�=�&*ikB�z�5T��7T��Y�m3�ׅ���ԭMsTpV�.qV�l��,e�fK�=�j�e�V�5��av�����e�i��-5gҶ�C ��0�Ъ�
1��94����gT�1f:4[,��7h�����e�-X1�Mխ[�f<��jL�� B��   �&'OZ<�k�,�Q�Sj�����Y�,OR붰�(�[d����^�VR�CY�̥2ĽIU*ֵU�j�mT�Sm�;b�̖�"����9��x��0!?��%|��>08a�(td�p��f�j��,rK���S��o��Si��2lY�z�U����ac��V�k��a��G��]�:|�i>6d>bj<�G��ǥ�*�:t�?��u"��,��N�S��\�>�d������R��)����9���i$��K%GK8��4��͛�aIVYf�3�.'*��Y�u���N�O��d�Q�h�gj��&JH��B��nY�E������Qg�G��n4]:<�W$����7��IЛ:��	5���������C���]�GT�OAy0�8�d�G�]��Ne��bn�(�o��é�:�����\��ܶ��<�Φn�soNtK*�Ŵ�����j�4=�;{#�ZLݧ*A��N�}~��$���3yԞ
R:٦�̖93������<S���W5)QE��9\{V2oP7IE��S�����h��Sq�0���Z;�g#lb4h���%���[D�.�Ud��,j򾆱��v�������IO��8�o_r�>'���7��x���1t���9���Iڝ�]�z�I����nF��Y�Pv����#���I�4v7�������U�J��IK�,�Nk�v;��:���ۛnmdM�̌��2떦ͽ-Q���8��jT��qq),����ū7D��D��ڮ`g�G���T���*�D�嗟)��5mY#�2d��МGSS�ް�dʔ�i����Ӭ���I<�*H��M�]��BCl��