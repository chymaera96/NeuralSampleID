BZh91AY&SY>�]� �_�Py���������`�}�@ �azy P
Ґ������ 2hh2�4 ��& �4d40	�10��D�F!�4� � h5?U@4  4      �H�M?Rz�����@   �$!4Ȟ�'��L�m�=G�f���m�D��H���'�?RГ`��!� )!X�`Q(E $B�(�����Ԅ�Q3T!����'�_esʷ���e�LI�yt�N�X���YS(ⳮ���'�S���Q�U�Z*`��I��>gR��P�%K�J\���t���S���N�I]�4�	��ٲ��lђ�̦�R�QͿ~˰˛��^���U𩜴#:��HI���3M���# ��h��$��m�Z�$G2k2S�j`���ۥ+g)H���~��㒟%17P�}}�GB������*�pḥ2�ӏIW��yHe���j	9��<�=�1wX��DD��#�aDƱ���p�-rK!-��;�j#���2���C�NjMdp)J�CE�՜b��X���ʺ�:��,��=e�u}j�J��JM��.l㉌
;�d���"ZP1FTr�6�',��{�8����C\���^�/��n9�IY4Z�a�&���C���YZK8S6-�b����t�a�@1ܘ����zֵ$Ѷp'�(�5�֝�}VhOl���J��5:���8�>j�8Y���MK�N��;�Z��,QT:M�*�{ـ��[3��ح�3��|X��:��n*K��3kJ�U�Vj����4�Ԓ����!�    �Lbp��Ď��7��g\���SĥJiu���� �I����+� �5CP���t��2����J�	�$$$$+�0Ɉ"&&�$R�#������(!��t�&KYt���Nʂ�D��Fړf��{k���N�='Ђ�5���uAM��وK�$YP�ۚ])����ѷXښ�)�d�6�N�����v����k����s�${�{׵Ų8:� 9P� ���!���mI��0�d�@R�p�S�$3E �t��B��d'�$d���}*R�L�gUBqE�䦒kR�	�{�U-->37�aP���Y���s}S%6Լ��G��W���i9(�A�u�^)��"Y��))��4�������ƶ�Zw�'��L��6���Vpd�Q�<L7'���ҥ9����Te"���a����{�(T�5N�,��z���O��䘔�]�I�� �a�
[�b]]A������d��'i����f�Ƥ�b�Y-���aN���&�&��G/"|�F���:g\H�='�
:��3y�'r�H�e&ǡ,ogSY�H��!�9�	�+�����r��o��-M�H6���/!�?2���0�c
�Yib�{���#2lLF�;���LL%޶�Z%Ԛ��Ri2�5;�ơ+��$a7�; �Y��[E(�EG	0��g��-8%�9y�u��oNC�w'cZ�'T��Xx<���j���O*U��Q#��H���tC�h��6��:�h�n�FR�*`*vG
^YV��g���t���f�&��Q5�l�.�3.�Z���f���s�8�3VR$ɸ�T���K�!�Q���	a�R�Sw��s0�4w���I�YS�pTJ	���/<Ƀ�j�D�?�l�3kPNu���`�v��L�H�LgF����S�Ȓ�l�����"�(H^�π