BZh91AY&SY���� _�Py���������`� �     � �`�2��j4I��� �     ����P � h   `�1 �&	�!��L��`�1 �&	�!��L����I��a4M0�2
z�Q����~�55=�7�
𐖐�B4����i	K|�O�Q�D��/
,�?U��I/�R#�f�ee����/�qU�GՌ�]<՟��<�,�o��-L0�����_��
z�z������(��Ye}m{���f���T�Oa^+3��s3m��K��:�28�M�p�ٜ��91Y1V�V���f5ɢϰN�d��v�#d��ϻ�xpp�Y���
����w)�Q��m6���Җ���/{�������j|K��6�ޣ|)/*���g}7��g�䓂��g�����&��e��S5��Z�)Ó��f%�b��`Yh �AmAh%�JPRTL�	`��ɺ��ڛ�}z�����{^i�pŮ�}Ta!���o-�M�4-. �F�-��SP��[�beQ��[��i��	�x���)U�UUUUUUIP����oz���>�l���YeQg�0��c(����n��J�[�j�Z�P_J�K��X�m�S,�e�U�T�*E)��se�2Z�Rp�:*R���l��uq��}s�Z��ow[���6��u��&����.ݵ5sw�9%�M/����Ѫlj�L��d��]U~�]���ɫS��|0�qG�96v�)�������ꑨ�*�Z�o}j{������)��g�o�:�/��|���O�8��R�E2y)#�,�6���c8�=���٣�aIVYf�3���VJ,޺�����O�����Xɠ�kWyQ����B��oY�E�������"����2>��Zg['���(�=FI��:�wE)�Mfo�FB���0�|>?.�B�h�%��^L#�=�|��ܘ��]��&�����v�tp���bn~ni�o[|w�SwFo$9���H��,[I���x�_��F��Gwle���r������{�ys7�I�#��6z��&pո8��8-#	\ԥE��R��=�:�$������/��)�40��aL,������r��14X�J���	w��ZQ��ji�5y����wC�{LI�$���H�_z�>�������n=�gd]#���k��[�w'Z��r��ȩ#�,=Kz4^Ȟx������b?'�rO��������@�1�QKĩ�<������gk�.��]����2&��F]2떦��3��qN�l��U�n.%%�w0yx�f�*G��w��s8��<��Hq�)�ة#���/>�dj�d�pɓ��IGF�'{�a�ɕ)�ѡ򧐧�e��e$nuG���"�(HWIH� 