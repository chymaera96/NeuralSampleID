BZh91AY&SY[��� ?߀Py���������`�z���   �0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`ba)�M�dz�i��F�    9�#� �&���0F&
� M# =LM0���FM��ړk��%��c3�����FR�4�������Gв����d��d��a�'����ߓû9%��xxSSHO��JQB�N����%��&2$��XHF�[��}E��+�g-.e2:��o2j޺�i���1�b�%�:�&-[�����u55s碙=D�ᕒDmi}��bw������s�Ud�D�
����w��S�d��].X!�`-t��eY*#�ұ�3U�&28C�K��s�lΔ{BK�01$�ħc�۩�j��	l^	�ƴ�y��[TM��$˼�NY"`�"��/���zo���-˖�K�r֫A|��5xͫ���(���Z�k9�N��S3��r750k7/���.&�sI�Hܚ�s�e:as����y�Н�Ÿ5�WD#�t�tUUUH`�&8����j�F��<TMe=��*.�ϒ�E�
-I"�~2N��#�)�X���΁5Ue��B�FK\Z�d�k�*�U"�֌����ح%i9��;U�m��U�������/�L����s=�Z�v/�������٭4qv8%ۙ�)�n/�mSEJbسj��U��mv��G�w[��`�ޓ���d������h<���E���F�֧�:_�`}�NH��K?vؔ�rw�b���G��7�~�JR�"��:i#�,�6Ƒ�C(��ie��'���(�qɜe�O�V*,ں����C��f(���Z�,Z[��1RE��b))�j�٬]���265E��7�bx��Z�g;q˂Q�y���$�M���4�L�������{���w��
�f�%��^L�^���˭0��]��&۱����99��w�M���<��m�ø�ɓ�'�8�K*�ų�GN���f��(���:��NNȟI�Q��<�N�),�W�,pe��a�ZI�W)QF˪���b�3r�m�����Ax?7�S$f`��`�-,T���L�2��a�X�J����]�3KB�4V-�b�����DW_��}�~*�S�pM�n_j�<O{{��?a��,苤u�i�u��pN��]��lS�t�H�3j3^&�'�*��{\N0>����37SsS�m�A�a��TR�*v��%.���8�Y�싨�gŵ�F֬I����$Ⱥ婳^��27�&��2V+Js����Q����ѓ�g�'��w���(�Y���r�7����T��~���Ϭ�����&,[���s.�M'c�a�ō)S�����S�e��E$ln&o�.�p� ����