BZh91AY&SYUrH� �_�Py���������`_z]�l*   �`�1 �&	�!��L�����2H5�      � �`�2��Jz�ʀ ��&�  �0L@0	�h�h`b`�!FCD�6�����4l�OSz�n��Ia�i#��%�0%-�Ib!Q��	�K�&d�#5H�U#5I��ғ���[�o�W��uw�L��,�o�OՆpY���ͬ%͊�FH�� �Cr��zM(��c!0��ےB��u��<��Cp�,I6,do湽��]��[�g-LSVx8�n�͢ϮI7C+I64���$�M=��n֛��j
P����.�:�����]9�O��r�[���LE��4�fΐ�%��v����B(����/��j�54� �e��X�ͱ�]�1���k����^�(/a099Ԃ!R��,aʈLg;ȍoQh�I]L�HAΐ��#8v�sCcIW�&oF���h%>�{�R`�M�д��	-�$�œ����ٱ��֘B��	�Ñ�%W+2��!q�WJ>L�D�t(2iG��)^S����LQrEUUT�I��ϋ[�,�Q⤛��,��,�(A
��v�aY�&$ɝ� y?A%�L\��\�	&J«&��
t�ArG`$Cl<CoBC2e�B���<o��{m�'��6S�t2v����]�����ΗmgxG���?1ǁ�4"�*P7�I}�������'�v�4�oz�8<�����ac�A��Ac�Fׂ�jqm|��E��Y���:.�Т�l���$ޯʟGR��H�bκH�E���#b���?U,��h��RE�Y�����J�M�]e�/{�qf�6�̔rv,f�ť��Q2RE��d))��4X�0�Y��[b,�(�����KA�������J8���t&��)�&���Q���y>����?_;��HjuId�y0�@�d�G�N�I�N%��bm�(�/��å�)�bkG򶭶;!����8�'Bʤ�m'��)�ؿCF�b�]qܴ���#5:]���O\���<�o'r���I��K�ᩬ9�C̜�!��*R��wU)N{�Z�M�Hm����Q����h��Si�0��!���r���,w%Ija����-�Ԭ��%�N���"�q��}�$��IO�Λ�M��]'���������3ܳ�]#��WYN�:rN�ܝ�jzN�I����ۑ���"yb�OX��~΄��976cluш��FJ���S�pRR�+Y�rηd]GN]��kZ�����#���Rf]r�׳�Pfot&��͒�K87���Q��ɽ���hh�<�����qh�f�*C���
�H~��/<#Sb�C��f�mjCz��k1;^E��&T�t�3�C��YO��yTT����2rE8P�UrH�