BZh91AY&SY� �߀Py���������`_ ��   0`��`ѐ��&��T�S'��&� b  a���b�LFCC �#O�H   �     0`��`ѐ��&��RB&FI��ba24��=F�F�&�n�+��d�$H���0%-�Y?�*%U*!uT���U�I.�f��f�L��ғ���\o���кb�⦏,[��-L0���۾?���y��;)�.QIX����Z���Jt�
����s3o]��{s��7�de�嚫��3�'���n͛�D2�H4g[�HtF.}��w��5R�UWs�]�;����)��w�K'2���aS���(�}g���Ie&�,���z�u37���U���q���M0�Ԭ�au�]
a�6T�ٴ��d�|��q�R���,�a�H��J��n��ad΍��cb�ڴ��ד'�i;c��	�2Ҟ�B>@  `���;ߓG�0Yڣ��<�)K(��X���k0��L�|���L���%�*����Z�ֵT���mT�Sm�cU�-Ei:�:ԥ�6��-��?��j�a�@�VCU0a�����5rv�8���^)���'�F���R�6,Ƀ�N���|-v��W�=nǩ��{��Gׁ�O?��Kl>�Q�S�AcЍ�*�bu7?��sE�ȳ�nS����J.v�k'М?W5)L"�:�#�,�56)�EGS8���ϓ7�(��ͤg���q��E��X�=��mY<
0�b�ӵ��x`�RS�3h�va޳1scj,�(��s#��h�t�xN|R���0ޞ�'Jl�:$�f�(�\�]������(Q���O9y0�0�2{c�N}��NE��bn�(�O��a��Ӽ����'��m��xM�ٺܛӕU%�i?g!N���Z4h{vx#��&nÍ"f�7k��=�J:�37�Iޥ#��m}ic�8j�aI!�N��%rR�Y�JS�Ǳc&�	�J.�MN��|_��h��Sq�0���h�3��F��h�c�*KS%ަ�h]F�ɩ�%�^'��"�9ǭ�1'�T��S�p��}ˤ�{���=����,ꋤvi�u��qN��]��lS�u�H��G��.�D��T�`�q0��_��>f�{i�n�a�b:�QKĩ�;�������g��Q�.߃sb�ͬ��#���4̺婳oSVg��٩L�N���;<<�t�y�{��`g�G���T����H��O,��:�VՒ92d����]ژ����*R9&3�C�N��E��x�T����?���)��M(