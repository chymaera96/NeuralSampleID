BZh91AY&SY �_ _�Py���������`� {    �& �4d40	�10�G��i��  �  4  0`��`ѐ��&��T�UL�  @     ��b�LFCC �#I&��b L&�4hSj=h�I�]�K�F�?��,���K'�Q�D��H��,�?%���\�j��Fj�L��ғ���\Uo{���L�ǝ4x�Ybߟ�ja��v����ৣ~�z5+%�(��*��r�%2S���N~��3��s3v�7���]vS}U��nY�F��SF�Y�����y��y��g�H��I$5��rC�j��s������Vi��
�����v)�Q��S����iI��T���M=s���3)݅����Y�%'Y_N���p��ѹv+����Lhe�F�����M�3�j�f��V-,aK6T�Z/����s,bj�F���m����ٚ�̛����x�w�]�-�;kM�6����8P��a�#@Hb���hH�M�mB��2�PZl�n}5&-)��!4  IB�OX�6Ϣ0Yڣ�ҟAJT��?E��]v�0��-*5�T�R����kUI>[�хiQ�jd�V��LMgI��R�Q��6]�%�ȡ�'�O�(�I��������?ݮ���t�>��j~=,�ϓW����ݵ5sv�9%�/�_��T��R�7,Ƀ�N�����v��W&�=ǩ�á�����y����a��ЍG�C�Acҍ�2���o~I��u���Y�7�t���Qs�H��O�8�~ε)L"�;ԑ�O�H��é�}��Ygţ�aIVYf�3�y\NUY(�z����L�F�'}��KZ�Jv�%Ix �RS�3h�va�Y����,�|�9���A���d�|����aПd��7u�Nk3}�2?gq���C���t��rY>��aq�d�#�N��ħ2��7ݔG7��a��i�17?4񷭾;O����9��"ʤ�m'��)�l�KF�j���{֓7aʁ��n��zOl����f�<*R;��g�,rg[�)#��yS���W5)QE���9\{V2�
�7�E�˩�^��S4ha��Ye������9�m�,xR��0�]�h���j����5x�SX���;������IO#�q��_z�>g�����n<��gT]#���k��K�v'J��sr�A�T��,<�;z4\k"x�ǴvF�����h������U�J�ӹIK�,�Nk�wݱuyv��۔olț�;Yu�e�-M�u5�\��tL�-igK��Ie�-Y�f��G��w��s8��<L�R�8����T�G�iy�0uF��H�2d�l�G[S�ܰ�dʔ�i����S�Sʲ�O��7:	����"�(H^
/�