BZh91AY&SY�"�� _�Py���������`�T@�@   ��b�LFCC �#��b�LFCC �#��b�LFCC �#	M������h�@ �& �4d40	�10T����&��f���SF���=���qv�KHL�H���i	K|�O��
�UJ$^YR~K�W�$�C5H�M#5+,4����V�[��1�������'���-���S(ⳲF�<<(�n�PD2#S��ַoސ�����gs9�����sSr�'EU���.\��rm�"OJz8�E�	ʅG;�M��d��^��bx�Z���wnp�Vi��UU������(�î��Ud��6�Wa3����d�ZY^�����>p�H.0��d����$d��i��&��D#�4�
^���k&�U6�q���3�zP������ǉ���{���h��\�
S�#*��B���T�W
t1X���u���w�E�*A��8�F"��f�Y4��gv���	B��$������Yi�s�mxF;|�6Jx��T]E��.�c�F%E�|�e$)��*`�I��'6�̓'wI��0�$��!A��	��LCh<�q!&d ��"��x�?���5�V$a�d�6��Ó�A|"�Ӧ��2��9Of��R�`,&DˎL�n�%��x.X�����sx=8t7�����<�y>vt<�5"��E���F�ҧԝM��0z✑a���K���\�>�d��z���)�S!g��8���V�MQL���R�?Fo��$QYe�H�8w��*�Qf��/�:�>�ř%l��Y��-�Y2RE�82��j�,]��w,�\�؋;�>O,���i��Y���9pJ:�9�B{d�)����&��ܣ!s�v�z^�~��H�R4r���^L#�;�=���.i�N%��bm�(�/��ÓtrN�[�qO+j�c���3x��МjE�Ib�O��S��~�����޴���*jrvC��=�J<O)�̤�R��f�t���55�RF��M�H�W)QF��S�Ǳc)Ф�l�];�E��>3F�����,Q?����r6F#F��RZ�a.�4KB�5+&�Hd���}mQψ�[�bO�%>��GB�WI�>����}泽�Y�H�y��S��9�J�nֵ<��Ia��6�E�D��T���C���	�4u�Slr��U�J���IK�,�G�:ݑu���[Z�mldMy���&e�-M{:�����7�D�U2:[��K(�������44T�3z�sR�q8�y��Ho���ԩ#�O�^}&��زGd����F��ɨ��v�>92�#�c:4>��Yi'�EI����ܑN$2Ȯj�