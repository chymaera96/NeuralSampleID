BZh91AY&SYD�Ԕ �߀Py���������`� �    `�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L����  @     �0L@0	�h�h`b`� �CD�L�&��4zOMM6��$���H̐�G�?E�����d��0��T�E�ʓ�^����"=t��f�i<�J��������iM^VX���-L0�����������}h��)b�JOMtT�:T�xx�V�k*�5�v��hv������pX����c��z�.[4R��l�M4٫W�#�lI���$:#rx�eϷ�q��ԭi)B����.��|Tnaꮵ���g:L3�3|3'"�T�K֍h��R����[��ҽ�m�qN&T�)ek�q��u8Qzm[�8��>^G̝6[%�У��S.��|欬��սdҪ�95h�e��s�&wi������5�_�Y�����l�Z������
�kv�՞9޾.�W_�L���8*��h�/��Re��!A   	��i�X����w��*M�}��)u~�]v���,V�}IU>9�ۙ�U�j�4�%Jlf׵�ke�˴��v��"��F��o]�+A���N��ʊQ~���k��k���^{���C�7��u2��-����]�}6sw�:R�-o��כ�d�l�L�,���UU��Z�Ŏ���=���Ë��GK{��'��'�����*����X�#��S�N��=�N�X|?��v<�Ԣ�|��I�Ȝ�?Wb��L�;i#�,��ܢ^m#��R�>k
H���ƚI�r:j����^�u����f(�(���+�Q�$]�"��pY�U���"�����Q�y�O��A���e�;:R���a�=�N��إ:$�h��d\�^������(T5vId�Ʉz���?�vw&%9�i%����s}^#�Dv'����\����<f�Ǝ�9��:��Ib����S�޿SV�O�Gw�=�I���$�N�|����v�ƏB�ȥ#��ozR�KHl�aI!�N����2���U)N���c.*�8IE�ϱ�^{�SDja��Ye�G�Z<M$4��1�X�%Ija���j���l��5�+<���Ews�{I�?�����)�+�]'��������;�Y�H�=��)��N��]��nS�;U$z�;���W�i�Pw>��'I�0~��O�����}.�#�U�J��IK�,��k�x��u���87(���7d�d�bh]r�ݿ����)�8�ee��NNE%�w0x�6hꚚ��%�{e�"sj�}����S�֩��<���q�z���.-�aк;����,ґ�1���v�󬴓ʢ���$���ܑN$#�% 