BZh91AY&SYf��� �߀Py���������`� y�    �`�1 �&	�!��L��`�1 �&	�!��L���{MLS �2    ��%=@2h ɦ!�i� �0L@0	�h�h`b`�!�44�MLh
h��G�6�~��	��$����,��F��".(���G��UZK��R#�H�RI��Rx��U�V����vׇ*jՅ�-�|��Q�e����h�ܚ�Q�,QINZ�}m����N�����+�f��e37�c��f���o�X����S6��igs����n��̙)�.�'�H�֒Hoe��$9b��MW=��]򪰙�P���|�xN�>�5a8Y=\m�s�y:�Ύ��)���`�G{�-�r������m$UR]K�U�S�-[��V��7�乿�~3ٓ;f�-���K�7��.Î*�[r�*Z�e���Li}�R��u(�	a�ҹa�6�N�#h���J7wzP�SP�Z��Ѧu�zѱTΓ8�WF�P�n�2�Mʭ B�   �-=��7<тεU�<�u�T]E�5�.�f��,V�ծxBi�3�)(T���(T)I���ww��l���cҦ˳d�(iI��
t(R��m��{+��k���N;zyܯta�?�;'��j���U۶��.��2]���Os��}4j��S&�0v)�U_/���X��jù���p��9�;�"y}l>�yQ��~qh,w#{�Sҝ��0z��(����k�(��$}�'Ԝ?gJ��L���H�'Ѡ��KD��g��Ygɛ�(��ͤg��9�VJ,޺���gC'��fIG}�R�X�YI��,�A�IL7�Ѣ��Y�j���͑giG��Q��t,�d�<�GA�0�Ol��7t�NY5���2?ga�������(R4t�d���'�?T��LJq.�K}�Dqz{�.X�N�s�qOz����Y�Ë�8�,�K�~�"����hѡ�Q�ߏ�i3u���u�q�Q�x��E'j���4��K��q�$r���9VF��J�7]T�9�=kNED������/��)�40��aL,��H�KG}��r6�F�;R��0�]�h���j����5x_sX���:���1'�T��c�8Hr/�t�S�������x���t���8����d�Nu�N��<�yRG�����q��⊨:���9�{�9��h�����ʌ*�^%N�ؤ��V��;������7�dM�l��S2떦���d���5T��pp),������7<��H�8.��\��'�7ܩU9]
�H�헟i��5l�G�'#f��]-LN�b��*R8�3�C�N�O�I<**H��k�]��BA�S�t