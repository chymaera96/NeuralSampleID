BZh91AY&SYm�� �_�Py���������`?H��ʀ   `�1 �&	�!��L���� BSOQ� �    � �`�2��j~�@  4      9�#� �&���0F&
� A224M4��Ѧ���4z4�M7�6`%v"Kb9��D�J[�d��0TJ�T��QeI�/U_�IrFJ��FJ��a�'w��*ߋ��4.����hɂ����S
8,����֧�9��˔RS��Z���M�L�u;;*�����Y��2�t��2km]v�a�X���
�;���&�EG���S=�,��Nhm��#&�U�hԞd�s���w��VI�R�UWc�]�9)�Q��Bf�p�vn �򢬗*&��^���n+��	R�C�q�M�En�ua� ���ǩ�3��Z�a����v�����C ���R�-$�){n��3[�s^Hʅ"��Wt�/��n��)wj��j��(�M��yjY�X���ޙ���b�%ǞH�\��h؊�K�=S�ђ-5B+C&4 ��F�b�����fe�X���V�MYDe�����H���|bň�aE�t.h2�m� ��  �$�M2�I6�ڞ����G�����,��Y�,�(d� q�Ň
��Z��&XwR������U�+0�ɝ�3	Mta=�K��ZJ�9��']J����J巍�z��~{|ǁ�2�'��\�~�%ڵ�GYcz]���s��x��5�*S���;窯���j,toh��r{^�[��F��S�=?�<�>�zP�y��Z�l}J{����&���g���qv�R��rG����S�qR���Y�Id�jixt2���K,�2}��Ec�L�,����U��6.�x)���kY:�`�,Y�N��b�"�4�J`س&k`�j̅�Mh�����1<�ah3U��^c������6��IΚ��Ni4�>*1?Wa���C�m�qB���K'���#�w�|#��I��줱6]�G�����S��j~	�ض��<Ʈ,�!��8RU%�g?gNֵ�ٳf{�rꏒ�d�o�)��Y�Q��2x);T�t�MoJX��5)#���̲%pR�j��Jo���bڤ��(�w�t������46)��,T��Z:�He#\a�X�J����]�f���h�Z�+<ﱤEr�9���I�U$���7H�WغO#�n|�j;��t�G���s��$�]��ԧ��T��,;���p�D9=�o0��������{[#�lG20U�J���IK�,��u:��8���ljQ���5bu�1�\�5k�h��rmd�k*��nn),��͹�'<��Hx7.��\�e�7���T��%9�
�H~��KϨ���H��mkf�2����u�8��#�a��:t��Yi'�EI�I����"�(H6��O�