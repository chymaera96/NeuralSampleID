BZh91AY&SY,oD 
_�Py���������`zAAҚ   �& �4d40	�10�6��D        s F	�0M`�L$$&�M(jd= 6��  ���b�LFCC �#I&����F��LSG�Q�='����I�ஔb$�G�>� ���r�XhM��%@&i~�6���L�"=T��$�l�Γ����*�7oVh�'ey|���u�-�>�R�޳���C<��ed�H\e����7&Z4��X`fv��3��������GR�9��.7:�"�/�s7YýRr�Ũ���	s�����$���$�5�A�7h�Py�>�t��UUt���<i]�[��9��`�{����vcʼf����>ୋ{ƹ���)l04�'�5[NYO�[o7Y�,�իZ[�^���:��r8t\�Y�.	��P[����ӫSKX"�؜L]a�81�@˵�����<�!AA�����"3J��b��b���A� �2�IXk7�j��mE�����Y�eR/*m�}Bֆn�3L��sY�Fo+0a&Ex[P���$$�>�5af�	f�����H�*�n��z���=0]ǌlc���m��m�0"�g�py`��0�Tԧ��(��>�I��]u�D��>�/�����mUVѻS�KZ��#(dbtlJi4��ȍ!����r�"��݋�����I�8b֊����%g᝻5��9>X�?�s��|�:����Xژ8������m	�ЩLZVb�ҧ%U}~V���˵�w{��ﻉ��Z�����I�a�CΉ�v(O�-�J5��~	�����|Sz,>���X��ou��G�L^$ة�oR��)����7"�����9YG��K,��~+�"����Y	��m��E��,a�r�yZ�Nw�Y�X�ZWAHb��:��RR�k3f���.�Y���ԋ:�<I��&��f�9���R�S�]Ğ�'"iޥ8��2|b0>��S���v9
D;K'��K��v�{����	yM���5��#s��.����^i|[��ֶ��:�;�9���MԉeRX�s�n�ja�͛3أ�<|֓'m�M�>��$���2w):Ԥs2MO:X��K�#��;S�dK�nR�Y�J�m�{1q)$k���3����S$f]��]K���H��h�e!��Qx͚�ZT���L�ih`�B�h3�ǵ�"�n�z����IO+jl�q0��'��l{����v�9c�t��e9S�r0pt���9�$z��sZ3`&��Pp{6����ͩ�f�q5�����U�%N�Ҥ�+A��g;�0Q���[J�mLI��������ji���&F��؜L��U�9
K(�ձ���ff�N���C�(���=�����R)�O4�y�����d��b������7�����,iHܗʌϥ9�v����EI\D���ܑN$�� 