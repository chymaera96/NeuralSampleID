BZh91AY&SYYX> �߀Py���������`�      �0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`b`� �#H��4ɂ#�2z�I�L����ሕ�$�I�5����i&��K'�(¢UR�^(������$�"=��I�,5����W%[�y��d�f�SW���-�?U��tY�w����O_)ΦT�E%=t�;1R�xxU)��W�f�W4�M�8�]vg
�9r�L�m9=��)��c���l��OiP�d�m6��Tj�d�s������D�)B����.��|�naڭ>μ����SE�1��k>z�D��
Y_?��F���U�S�͖�ˌ��%r+S�+_u3�N�YY�r�gV���8CJx�h�\]�I�:�ʱئ�LT�}5�W��.�8j�l�eu�φ4�fv��n�t�]�[�����x��U)JR�����������Otx��s�w���7�}G��*]E���]��0����7ԕS�l^�V���r�dқ4h�UZY����"��E罽v��J�:��;��&�����/�k���^���n��o���e���??��v�l��,sK���S�^����y��2ܳ,
u�W��Z�Ŏ�m�{��k߇$���{��'��'���C�&�Ψ�"�X�#��Sޝ��0|"����K?ӄS���~�;䏲2������R��)�g��:"��km��#��R�?V���$QY΍cM#��s�ʋ8.�x��e�7�̣�͊]b��z̪H��E%0�F�af+477�����2|�h5U�l��o4����qO�I֛�T�T�M�����������NN�B���%��/&��_t���LJt.�K�و���L;]Qڞ&&��螇�Gy�7v�y#��t�,�K���-���j���wyc�-&��D�)����}rJ<�A�Ԥ�R��h�޴�ͤ6n0�����R�a+����u�JS��ֱ��H�$�����/��)�50��aL,���Z<�$4��1�X�J���	w��ZQ����2����DWwA��ğ��%>�4�W�O���>����K�Y�H�=S��)���ֻ��ܧ�y${KK���W��ODUA���ts1?��9����qo=��#�U�J��IK�,����y]�u�����pod��w�g�4.�jn���499�$�4VV��rr),����ɳG\��Rz��~�04�ѫ���*C��N�b�T��>�y��;#f��:FYqok'R��lbw��Y�#�cJ5>4�����΢���$����H�
!��