BZh91AY&SY��P� ߀Py���������`� @    9�#� �&���0F&"��z�*z�P      b�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`b`�!&#)��0����mG��6�v���	��$��Y	K|VO��
�UJ�YR~K�W�$��"=��$�Ya�'��|W��ߚ.����6l,�o��Z�aGJλ��E<��#
X����έ��*d�����nV��ܻ^w3��5��]v��jmX�ߝ�.����p�viX���S%8���D���$�͌������6.}_�]�����QJU]��w��S�c���Y�^�\u��t�^i�VFJ��+<���i�ul��Ȳi^��Y�tITd��K��W�i?�RB��,߲��3ц��v8�F���Δ�m�,��Cu%ZЫ�;�&Yk�����yR���/X�����iԲ�%2�jb�HBbHh���0C&�@����J�<nmkk��,�6��o����z�JR�[�UUUUUT�,������#��>JmS�<�YE�Y���.�kae(m�*�����V�������2��R�њ�r��ѵR)M�e=M��d�6Ro}�Ϊ���6�^覆�����t�����Fi���N-^���f�j��,qK�^)�}����UJdس&�:j���-v��W�=nǱ�á��qmu�������!�F�ġ�E���F�ORu7?$��sE��Y��
t��߹E��#�>D����Ja�YऎH�|U�FŇS8�y�e��G�(��ͤg��j�Qf��/�:�>vՓ�ر�AbݥI��,���IL7,Ѣ��Y�z��͍�������G�n-�����s�uc���:Sg5)�Mfo�FB���0�=����"�#G9,�Ay0�(�{c�N}��NE��bn�(�OWY�6���&���3rۣ��9�x'Br�YT�-���;�W�hѡ�Q����f�8�3S��}~s�$�����U'z��4��%�,�a�$o1oYJr)(�uR��q�X�Ф�t�]<z�E��>3F���)��X��h�g!����Ѣ�zT��K�-к�U�SA�Ư�k]��`��&$�
�S�qN�]'��8=���67ֳ�.��yg%�S��;�wc��O��*H�7��.5�>h�����������:����9��ތ*�^%N�ܤ��V�%�:ݱu����nmdM�����e�-M�z���)�:��U��.%�v0xx5f�)W�[U��rh�3}*���S{�R)�y%�������d�����G6�'k�a��ʔ�I����S�SƲ�O��6:	����"�(HW(~�