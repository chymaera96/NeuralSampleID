BZh91AY&SY̬�� _�Py���������`�zQA�T�   �0L@0	�h�h`bc�0L@0	�h�h`ba�z&�=OSj       ��"�M@ h@    9�#� �&���0F&
�  # M jh���zOMM6�n]��1�g#�?E����,G؅C*!P$b=J+�*Dz�|�L�$�Ya�'���\Uo���拧��ʙ�LX�ς����K;n����^����ԅbPHi]m)3���P�n��>���uu��dp�����u�����\�n6�ќαf�.�a�����Î-�ީ#|2��F�������>���s���E�"��|h�h��.%�g��(st��s-3���1]YS\�g��xsk��%%�[��m��)�͔_z�¦>����2c�έ%7*�4��YɊ��c���L�JJ�j��^���lf{��u���9���ʖ¯s�8g�[%�V��FA@���`������3q�j3tbK�NǶ�罣[5a7]lf��±��{��w�"". ���������a�;T}U%=��*]E��������D$Io��H��f
6������֪�hʙ_�v,��ʔ�%�b�R�(�{f�h1(kI�����J6�q�	HS�n4$��Y�e��������������M���)v�w�}����͢l4T�-Vb��S���]�c��F[��{pnp��8�:�d����}��A�P���X��kʧ�:[_�`{b��X|�?v�N�7{�(��$}�Ԝ?W5)LLE�T��E���m"*,�����>l�k$QX�8�!�p8�b�ͫ�^�t�x�c(�cb�X�b�;K�H��B��6�͚��,�޴�\ձw�})��KA��蘼>)Q�y���$�My�M�i2|b.~�������:
FnrY=��a�b���N}���"줱6݌G'���;9�y���9'��m��xy�u����U%�g?g!N����f{�vu�ⴙ;4���I�Q��<�N�)L�d�,��S$o0��7���)J�5��Jq��,c7*$�%O&�Ix>O�L���n�)��,T��u��ț#͚�zT���[4�.�Eb��b����DWg!�=�Y���RJx�S��ںO��8=��5<��Θ�Ga朗YN��N�ݎ�z�I����6�5ƒ'�*��{�`�`0>��qO��������0�0���U�J�ӹIK�,�K�u�b�9�����Q���5��bc�2.�Z���h288��2b��Y����Q���pf��<�)p]�h���'&o'ةU7�U"����^yL�ѱd�C-͌ѽtsha;]��4�rL2�3�N��E��xTT��q3�w$S�	�ȝ@