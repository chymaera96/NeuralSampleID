BZh91AY&SYm��z $߀Py���������`� u�    0`��`ѐ��&��T���4�PF�@ �4@  ���&��       S�R   4     �& �4d40	�10T��i4Ѡ&��a0�SG�4�=����!]�Г)���|ֈ����d��0��T��yYR~k�W�$���R#�f�Ya�'پ�U�;{��t�)�����>KS(Ⳳ��z��f����yrY��J���/˞4͕K���T�?��ͺ��fi�cy�����7,d^�h���t���pli�e�T�-��a���|5���l�\�jxj���mnެ�d�P���|�xN�>�6��sU�顉QT�9�|�S61�ƅ������]�6R�j4R����'n�4��㩐B�)aQP�)!��L�$��d�V[�U�Z8�Y�k74ɳ���h�*���-SJ5*L�-Mme*Lf��a��h�PJX�d����1'��kTkp���ʍ��]���yh�{o�s��EF9FKU�ԙiO@�!!�  0cI�Y���^X�gb���j���YeQg�c�Յ�K(�Y_�u镊�B�k�2�f��1�����K�Z���lYy��U"�֌硪�-E����;hUJQ��]W��\����?ݳN:�9����Z�fO����z����M�.����������ѱ56*S&ՙ0v��U_/���X������y�l9��G���<��}l?y"lH���X�#s�SМ���0zb����)��w?b���G�#'Ԝ����JS�BΚH�'�[[�J
�vq��R�>L޶�Ee�m#<�w�NY(�r���s�}�Ve
:�k��gaP�Ix ����h�b�,ùfb�֨�����L���ņ�E�̞��Q�y9�$�M�
S|�&or�����a�=���+�P��:$�yKɄx�{'�?T��LJq.�Ku�Dqz:�:�;�M�{�x���������#��N4K*�Ŵ����sU��4hz�u�G�i3u�*A����1�Q���jN�),�W�,pg�����;�z�0��JTQ��)��Ա��P7IEӿa�^��S4ha��aL,��Q?����C9�#F��RZ�a.�KB�6+&�I,lx_{dEu�r=/9�?�����#�}ˤ���+��=�ӽ�Y�H�<s��)���i̻��ڧ��T���r4^F��Pu�C�G0~���CGS���n���1хQKĩ�;T�����q\���Qїg���F欉�#���Bf]r�ۯ;d��W�NFj�KZ�g+�����+c74�4Q<nU�����qh�}�����Ω�O�^}�x��d�22d�j�&����bv;V<�R��1�t��Yi'�EI\����ܑN$}o�