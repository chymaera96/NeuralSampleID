BZh91AY&SYq� �_�Py���������`� �    �z�mOQ�h&@��4� j ��        9�#� �&���0F&���        `�1 �&	�!��L���� L��4OS�#&��44zM���M�ۄ��Ȍ�H�g�`J[�d��0��T�Eҋ*O���-Uh]j��Fj�2��JN��TW����]/W�l�Yb���0u�W|-�������f
)+V���jvvR���+�g-w3��k����ˮ�ر�͝�.��K|�ozYiv�gn��T��S=Q��hHh�[pHsF��&�ϳ�j�ݽY���
�����u��[)�_]��Rm7/�!�%K��in\K|cM�؂�MJ�Q�T6S�ml^b���}	�\�Z�ʬV{�ϡR�-F�_&y�V����+^��V����V��.(0hp	jC�AM�r�0��R�
R��40�m�*2����%
2BC���3 %��!A  	�cI�YLmuOע0YN�X���OAJifE+
X��ZOR�0�L�Qy��i��k�V2��5-MX�l�_FV2��z�Rغ�R)M�}LMk�d�(j��Sz���T�BR)�c
���=���F1���k�����H>�ײ��]��	v旊}����Rl5*S&��0v��U_/���X������z��77������y��|�>�yơ�R~qh,zQ����'Ck�L\S�,>E��jS�����.vI���&�O��JS�BΚH�'�A�EʅGC8�}4�ϓ7�(��ͤg�w��Qf��/�t2}�'S�c&�b�v2RE�H2��j�,]��w,�\�؋;�<^i��M���*Y���9pJ:9���I9�_%)�&��ޣ!s�v�z��~?��8�CG),���a����r�LJq.�Km�Dq}]F���;�Mo��<ͫm���k��Ҝ[��*�Ŵ����sb��4=�:���ZL�g
I3S��=���$���3x);��t�M�:X����)#��;әa��*UUY�J�p��,dܢM�Qt���/��)�40�m0�Yb��V��r���,w%Ija����-�Ԭ��%�O+��]|GZ}oY�?����|�ںO����ͣ�5��zΈ�GY�8����	֜�ݭjz�I�ý�ڍMR'�*��{Zp0�>��pOGSsa�m�A�b9��QKĩ�;T�����q\���Q�.σkZ�����#���$̺婯gCRfopM鹚���k9���K(�`�ojf�(x7���.`g�G��ک�59�
�C�O�^}&��زGɓscA̺95��Շ�L�H�΍�:Jw���ʢ��m����ܑN$\F+@