BZh91AY&SY2�Q �_�Py���������`�z�T*�,    c�0L@0	�h�h`bc�0L@0	�h�h`ba)�&���= Ѡhh  &�
��Ѝ0H��0	�� �`�2��*H�hL�D�d4$�G� �	���M�لEu�$��Lb&rO��R�B`
+�(���PHId�2Kj��!y$d�I餙(���#:N����v�v�ҾIp[�O������<J�ZZQ�g]ߟ�V�֣�o���Y��X�E%o%�����$A��mB~q>���[=����9��L�\�9��˙&�a�c�I#q��i�V��J�et�5)J��RI�F�$��k�^&�1hS[�؟����ӏ-�ՠ�"�J����ș��Q��ʅ��g�	ơ\԰Θ�k*��ٲT��}�n328��1��ו���LHt ��<U�n��a�( ���<����70t4�:l���|Y�嶲)lW�=V���^rVn	�<F$Vza�n�d�j� �;�]��=�1Cj�Q�	^�ʲ�;5ٝ%A��&�jA\�6�4��{�0RX�� ��BC<�EŒ7�&؂�1����՜Н��50p_h1�q����EUUUTB��ROѩ�����=�e�j]��O���AI$�p@�ʹg.*�dT,���X�2T%�3$ʎ�;�N��ҲKD�����&-�f!ayqP%�$/I�q�dUbLT%��k��z��?<{���f�(>�C�p�����c(���7���%=ﻁ��Զ��4TS&�̘e9������L�S��=����񓝖��<>���C�I��*G�KI=$��)��1=rQ�$������s��oآ��"r����I�����JQ�)�,�O�ҋ��M��B��������>fOsP�qɜe��3yЪb��,`]�����],�vŇb���b�4�`��K��2E%1mY�2�v0w��]4kE��C��LS�F�5�,�b�N[ғ�zS�!ΚqR���2}�LR\���	�~�gw;�(TM�,�-K�<�����^$�S�vP�M�1�8�}F#�8��h�
S�w6-�:��N,�R8Q¢Y*�al����x���3ff{Tut��-�I���E8�)I쐣���O9Iڢ�Ɉ��K�CQ��I'1�;�̴��e)(к��7�{L[U�"���GB^#��ș��b`��,RO��t���&�0�٬v�I{���]�3����P�F%�O��"WW�#��H�EAN�zn$ھ��>�����4;�z�D�I:�4��s��R9�u:�)�r*I=%�{�ߴ��$i$���Z���<R:.21>��	���m���m��6$۹�IF;d�tY�rYZӒ�'d\��ϋi��ֶ)4�v1LzFE�KQ�׳����{�7���Tĵ�q7���N,&��#�f������Թ��C�����*wԣ��T����y��`tI�ֲI�Gݓ#���$ܺ940��b��bƔ�)�Tf���%<Ŗ��T�hړ�|�"�(Hg(�