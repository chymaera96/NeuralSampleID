BZh91AY&SYM� =߀Py���������`�@\MR    s F	�0M`�L4FJz�� � ��  0`��`ѐ��&��SԄ��&��=G� hh ��0`��`ѐ��&��RD&FF��z�6��MM�I��m&���bI�#9���H�J[�d��0TJ�T�.J,�?���\FJ�4�� ���<7vQ_��ߒK��7�I$'��JT���N��%�z�����*$%mn��j�]L���4�W��圵����[�n]vfŌM�\��u޶��X�l��^�*��6p�vO�m"#6�m���S̚�}��M]�hJP���~k��5<�j��T,鯪�u�Xƛ�,1�1Y���f��MR_\���4w{V�*f���I������4�u3�r֮�7c�����g̖4��"�.j&4u��II��$�!��q��.�D�� ���j���#�P�U)Nw���&e��@�,��1TڧI���)��
TI���4D��+���̶�5�$�g<�����p���UUUHB$��o9��*n��})K(��Z'��0`�e�k1����Vj������
Qi2�Q��i�+�b�s��ѱR)M�c>���X����F��#j����ܥ'O4�,?�X��C�K��ac��dq�r�3�dm7�����_ߋ�6���R��Y��N�����R�W��7��������zS����a�CԓA�Q?�=h����S������ȳ�m%:\��Ԣ�l���ț�?W%)LLE�t��O&�!zER��eo��Y�2}��Ec�L�,���p��E�WX�?��b��N�2�b�n��j��"�4
J`ڳ&k`�z̅�[gyG��1>D�Z�gK���(�=F��t����D�L���������C����"�$��K'�^L�^���4�S�vRX�n�#���0rtG$�0����6��;O1�&N�qnN4�ʤ�l���)�ؿK6l�j�}��V�'3��NN�{�g�IG[�d��;Ԥu�M�RX��50RGA�<�d�%qR�Y��J�q�XŹH6�E��3��ĦH�����LYb������C)#͚�zT���c4�.�Eb�̘�h󾶑ψ�O��0���IO��7��ںO����ͣ�5<��Qt�g�q]e:\�t���j��u�H�,<��f�4�=U7�s'`}����Fn������h�:����T��J]aehq\���Q�߃kU[�\N�&<�"떦�:�#{�oM̔�iN����9�<��2t��ԓ�޻��s�N,�vO�R�Jt:�"�~���Ϝ��H�LX�63Iк940��凖,iH�eFgƝe<ZI�QRF�����ܑN$pC�@