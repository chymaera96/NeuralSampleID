BZh91AY&SYf�s �߀Py���������`�E��   �& �4d40	�11�& �4d40	�10�OS��jz�!��bdM4���� %=Ji4� 1    F���b�LFCC �#I&� ��L&�4��P=&ji��p�Wt�#!���~kA����d��0TJ�R"�QeI��U_�IyJ��FJI1��:O������8]<�v���BI	��JP��Y&�G���������bZĨHb��g+b�.\Q2�A�����S#�u�����nX����3���)�qd�0���u,d���^����Đ�ٳ,	�;�b����qp�Y&�R�U�>
���&"�	��n�x���I��;/4`���d˯*��E�5.�{U}��٬������,uTE�$�YV����e/��qY]��o�>�Փy�����3n��n�&�]h�e����J�[m/X��]�-�z�Li�J�T�ݩuI�e<�20ſe�U�a/kޥ�?e�Vmr�}p�f�j���]��EUUUHb$�ۈ�_-��gj���YO���eK���X�uڔ)BD$m���2�2�^"���,�zZ�h��ٰ�Ŕ�-e�5T�SZ0�ƫ�b��5�����QJ6�k�)Cd�������>t�q���A�0�ڐ0���QP�h��,qK�3�S�^O�mSEJbسr�U�|mv��O��c�����>1ū��OG��K��h<���Acҍ�2���m~)��E9���,��d�C���\�>�1}	�S�sR���Y�I�d���ؼ:YG�饖~L�s$QX�8�)<\5X��j���t�}MVc(�cb�X����j��"��2���fL�.�f�������1>�m-j������(�=��t&�jS|�L��������{��><�C79,�Yy0G�x�{���>��S�vRX�n�#���`�����l|��ڶ��;͜�:��ܜ�U%�g?W!O��3f����돊�d�8Ԓd�7l��I�Q��<�O)L�W�,qe���)�h`��JTQ��)��ڱ�ܢM�Qt���/��)�30hm0S�X�e����R5�#6k	RZ�0K�l�к��C91X��}�"+����z�$�j�S�qNn_j�>����6����{�t��;<��t8�bt.�w6)��J�=E���ڌדI�Pv=��N&`~��qO������m�a�aт���T��J]aehr\���Q�ߋkb��X�f'ki�u�Sf�-$���tɊ��:
K(�`w�h��33T<���0D���d�U!���J�T?d�K�1��5Y#���nj��G6��ܰ��cJG$�*3>T�)��O"��677�rE8P�f�s