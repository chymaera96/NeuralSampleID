BZh91AY&SY�� �_�Py���������` �V�   9�#� �&���0F&�S�@      `�1 �&	�!��L����I�LѠ`#��#` 9�#� �&���0F&
��# M ��jhѣj2zOOT�i6�Ew$�@Ȇ�?3�Z&!)o��(¢UR���T���U�d��L�"=+#E"ge��O?ouqU�7�ˤ]1X�SG���-��0K;n��Z=
V�&kҰ����7]�=*wwU)��+ĳ�;��͝V8�\]��c#.,�+5�&Y�S޺��8ݣcֆ�e{����	�MK�g��Ŧ�f��(UUWs�Y�;�Q��S�}W�L��n�]ٮ���t>�L�wk{[&ؒ�K�e|^-K7�}��mW�7��{Q�fk�������.���f�͒뭛,۱�M��}-V����imVe��LaFT�G�+K[<��	i
���m@J� ��P�5øW
e41�<%��r|Rou�BI@  a�*{'{�5>��gj���%>����Y����la�Qb�4m՝�Z�,��GN��������T��ݔt3*Se�Kb�-Et���;�)C�kA�	��c�_���o�$d|,p��^�jrv�8�ۚ^)���'��I�ԩL��d�ܧEU|��Yc��Ss��=�np>ű��'��'��5���ǩ^u>��m~���s�a�,�e:��آ�l��̟2pT��ԥ0�d,ꤎR,�
��j"�K8�}T�ϓ7�(��ͤg��8j�Qf��/�:Y<��'Z�3�-�S���x��RS�3h�va޴�\�؋;�<I��MBΉ��s�'��r{��	����&��ޣ!s�wz��~�@�Q���O���G�y�=��S�bbS�vrX�n�#���0��Ӽ���ܓ�ڶ��<F�l�So%'*�*�Ŵ����{b�4=�;:��ZL݇�3S��{�G�IGS�f�);Ԥu3M�Җ8����
H�bd޴a+�����jR�n=�7*l�]<ڎ��|_��C��0�Yb��Z:��fM��Ѣ�zT��K��к�Jɨ�d���}mQ��vO��1'�%<�)�I�}����k���>�Y�{�t��;D��t8�bt.�w5��J�=e���mF��R'�*��{Gd�b`����<m͇��9�шތ*���S�w))u����g[�.��.߃kZ�����#���4̺�jk���388��3R�*�Ie�.L�ѨԨ���{R�q94xپ�Hp���ҩ�y�����H�2d���7��mF'k�a�*R9&3�C�N��e��x�T����?���)�(� 0