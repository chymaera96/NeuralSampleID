BZh91AY&SY&ݕ� _�Py���������`�*    s F	�0M`�L%4 ��Dd� �  4 0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��RD&LF�'��2d�Ѡ��dڛ"oRl`�v�,�1Dg#�|��	K��O��D��D���*O��U��.��R#�H�P1��:O�%nU��vc@�Kv�dT�����D� �������['����`��))7Yu2S���N���uis)�ײ��&�Z���b��kst�w�lj�Z�N�f��d�OT&�eh�ji~�	ю�S�4`{�ݭ�U�h�P���|�yN�>j5LN���Ǎ3N�GwV�F��t�P��(��������V+p�x���覌��D��?0�,�r���A���S��:�-��2�!f(ٜl�F���8�f"����1tf�&���`���L�}�Ιm*P$�Z�(K�D��6���˽<AUb�q&|�[ޙZ�wWK��Бq,�ϋ����!-D�I$�C!���8_���v(�SZ�����Y�ZG�$�G;&��f*���ҙ�ei��pzC��.$8��X�KXr*�ƵH�5ь���d�h1(k��$�L$�f�����y^/_�{oc��jx�����=����v�t���Xޗmgx���8�y�Mf��ũf,�:j���Z�E��0{\޷������y�������"��Acҍ��O�86>)��rE��Y�6"�.N��Qs�H��ě�?g%)LLE�T��O�SI%�(peo��Y�2{X)"����Y#���U��6.�xY���kY:�`�,[��v1Y"��2���fL�.�f�����gyG�嘞(�Z�gKq�zQ��6��IҚ�)N�4�=�1?gi���C��nt�Lܤ�zɂ<�����r�Jq.�Ke��q}}fN���S�qO+b�#��5rd�G��D��,[9���w���͛3أ�\�����H2S���I�Q��<�N�)L�[Ζ7���F
H�0��t,L�ҕY�JS}Ǳc�d�]<48����d���e�*'�Z:�He#\a�X�J����]�3KB�4V-ъƏ#�i\��h���	?�����tF��.���[�������g�G3�8���-��:Wsv�)�:�$z�����$O,UA��Ѽ�s�7������}M��6#�*�^%N�ڤ��V��:ݑu���65(��Ě�;��L��Z���h����6�V*��������l��:ffj'��w���(�Y���b�7x���O�>�y��#F��8�-�l�к940��Շ�4�qL2�3�QO��yT��������)�6�@