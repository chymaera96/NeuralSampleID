BZh91AY&SYkէ� *_�Py���������`���   s F	�0M`�L%4"T�����=CF�i��4d�	��s F	�0M`�L5?U   @     ��b�LFCC �#I&�	�����dLM54z��<�z��Ԛ�!]QГ������������]Q*�I#	YR}XUW�$�Hd��d��a�'o���U��]�D�n��J,v	pg�tI"C�0z�7>��m#>J���E%wԘ̬��S���No ��6���~��bLA�l���5�Q��i��9���'��AT�v��\Dlh�e�Hҝi����͚Zu+$�"�*�����⧊�-����kۄ/�S�Y���j��r*�P�R�\C���b��!�\�b�a�C���^�����J�n99~��*_'dmT\���ƔlD��V�
|��u"ڎ5�x�0$�.:�+��H,�H�"���[w'�j	$��J�p�>̗�&bH6"+Ud���^����z;�k+? �Li�:7V"��A�ԙiO@�!"   0cKOd���hw��:Ty)�S��*YE����dh�I@�ӷ�����"����Y1(.C�%�'wI�@R.<	RcBf� �w\��
P� �Bf�d6�D��x^1o����s���&���(�s==���:FGH8s��w�ۑ﹁�"��Q!������?3B���ci>q����OWȞV�=Q42�}b�X�F��O�9��T��pE��Y��ȧ+���(��=�1yj���JR�"�zHދ'���-R'3(�<)e��'޺�(�qɜe����uV*,��cI���jY:�L�b�*ºJ�U$Y�B��kY�5�Ywb̆��Y�Q���O)�ԋ9X����c�]�>NT��JrI�d���`}�E޷�?��(�Q3p���a%��;X���)yM���5��#{��.��	�^i|���ֶ��:�<9�olM�ʤ�l���)��Õ�6g�G��+I����)��#��{��s��N�'b��vI��K�CCIu$r�jr-�[ԥEiR�݀�,c6(���sA�}
d�˴˩u�X���h�e!��Qx͚�bT���L�ih`�B�h3��Ƈ��h��;�װ���RJz�jF��$�?���|�'kⳚ0H�wM�S��8�+SJ��:��Ya��kFl$h�<�U�q�������7'������5� �/����*uN�%0XYZ�:1������TkjbM8�,Lx&FSN�f�[�jl�*������%�q\�����33TN���C�(�ټ̞�Hm�S�̩�OL�zK�ѡ�d��1b���'#ph/:]KXґ�/��Js��Yi'�EH�M��|�ܑN$�i� 