BZh91AY&SY��c� �_�Py���������`�  
    5M5z��&�F@�i�� �h���b�LFCC �#��b�LFCC �#��b�LFCC �#��b�LFCC �#I �L&��4i1�#�i�&jjoRpĒ�`�������Z	K|�O�Q�D��"/%T����-Uh^A��G�H�I&l�֓�����>ZB�z��4h������
:�w]��ڽ�z���z�*\�����Zr�E2���Jv{��Y�K����YwR�7�d���Sܻ��y=̳�s}f�+�Wl����p��i��TnO:n^?w��s�5h�IJU^/�w��S�s)�V����N������Ě����j�:�����Sx���&�,��k��Z��:��]K�Z���})k��*о�r��*�T�M���z�μ+M4gss]���7��[n��f�b�سcZ���)�V�q-��k���vmfr�����6�ὣ�gٍ2�[���h�zp�ugw}o%R��*��UU*���*K-=�y?Ã�ܗS�V>j���������걲뷰ƹ]E�%�U)����f���S+�miT�j٫ŭf6Yv,�oT�S}[z�Z7R~��C�JT�*o޽�HQ)��Ic�T&@P ⨢"�&{�(�r��iw��}���|�l�͕)��`�S���O��n,vsl��w��~\�����Z{?|�?�=��z'��ǹ�>��p~i��tE��Y��$�[���\�>�2������)�S"�5$v���j,ܴ�RTv4���K,�?s
H���ƚI�r�EeE�X�?�v2�[�f(�Q��,�)੕$]�"��pY�U���%����g�G��L�98�j�g[/9ӚQ�{8��$�M��T�M��������}���ד�P�j�%��^L#�=,���)ӽ1)�]��'�����::��y����>��G��7th�I�❵*�ŵ���)�޿[V�O������I���RI��~��$����'���3D��%�m!�q�$u��:���j��n��Js��,e�Q'	(�zv;��|Jh�L68S,�H�������7�#V�IRZ�a.��KB�6V[ɕ�����"��G|�c�bO�%>�4��.��}�O��~&���vE�;�\�]e:�ӽ:�w�[���eIQa�z���m"}U{�;��bL���i�5w8����#�U�J�3�IK�,����;�u3��87(���7d�d�Dк婻ci499�$�њU����Ȥ���?&�sSUC���l���N֯CGک_5:���P�iꗞ�dl޲Gl�eŽ�:�GF�'��a��4�v�4�S�O1OJ�I=
*H��M_�.�p�!����