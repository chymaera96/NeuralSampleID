BZh91AY&SY�*� �߀Py���������`� ��   �0L@0	�h�h`ba�Oҟ��z  h  h4�  `�1 �&	�!��L������S�`�&�L�C M4h��0L@0	�h�h`b`�!#C$�Majhѡ�4z4�6�v	]�"�2!���~�$����d��0��T�!r�*O�z��d�j�U#5H�Ya�'gmoU��ɢ]2�t��ae�~%��pY�w��ѵO>�^zע�h��uV�K�%;{j�����Y�]��fͶ7��]vF匎}�,ɿ�b�L�,�_~u�Իɛ�C�֐��\��S�}��v�?2�MJP���~��G%>j60�tײ��ZNE�.ͅM=N����Oj��a&�*���c-�A��m��/S*�)�cw<�e�ؤs�6��n�+/�9�XYu˫&�0�l��V�igJ��U�מ�m��u,�B�[/��#8L	0���$6a-%�ƕ�,���s������JR��ܪ��������OQ���^��gb���T��,��Y�-]v���-*�^���mIU>v��/U{Z�2��)U.Rjfͣ�YL�6�E)��O[b�-E���䜔R��1�!=(��>��`�*����*�a��m5pv:�f��}����Ѫm5T�M�2`�S���_]����Շ���{0�o��t6�2y��},>�y�Q�Q�E���F�OZu7?$��qE�ȳ�n)���~�;$����&�O��JS�BκH��'ͤ6(�
L�����>L�c
H���6��g{y�U��7.�xY���mY<
0�X�݅���.������f�b�,ùfb���Y�Q�x�G��ZgK'��Дusd�I:Sg)�&�7�FB���0���~�B�G,���aa����8�LJp.�Ku�Dpz�\��;�M���<m�n���l���ps'
K*�Ŵ����sj�-4=�9x#�-&nGEf�a����%o�̤�R���6��c��5l0��s�Nu�	\�E.�U+��ڱ��H����ߡ�^��S4ha��Ye����r���,w%Ija����-��Y542X��}mb+���=F$�$��Л���]'��[�������gT]#��YN�BrN�ܝ��z�IQa��7#E�dOUA�������	�4xͧ��8���FE/�l�RR�+S��d]G�>͊76�&̎�F\S2떦ͽML��ޜ���iN����90xw�f�)<���W03�������C�NwR�R	嗞STjڲG&Nf։κ8�1;��L�H��΍�:�w���Ģ���bh���H�
\r@