BZh91AY&SYj�>� �_�Py���������`�zQUt@   9�#� �&���0F&���z@       `�1 �&	�!��L����&OT���=M �h   d � �`�2��*I4 ��24&�)������S�ޤ�t��ȌR��G�\J[�~�.0��X�P��,��Ib�R#�H�Q&6XgI���T����2'evޙ;WYb���.��:�}>y���6����G�c�L�d%�۵D���Y�fS#�E���65ҬbV��ʛ��og��7���]���#l5Z1�rCliOi`{��*���IJ�ӌ�������
���/W"��
R�к��L�S{�6zz�n���0���5�3�_V̎S+�l�e�Qfֵ��L��54�lߛ��Х��M+e{����5����c]I�Ɋ�Hd�&L�{�2 ��0:�n�� �Jk�N���i �-�E95�q_Ma�<�p�����OhN��(���UUT�(��'�38ap��!�8A�Q�T��Ō.\�
�#��\L�A}MLʨکj�d�����ѵC ��-;���fE@2l<�� �!��-c���մ��4��f׾.�O����w�>~�:����Xޘ63��{w�L�	��bdk(ȸm����V4�9��.��;��ln��ڝ/2y�$����j��AcЍo*���k~�s�qE�Գ�kJs8�r��#ؘ�	�S��)tSgE$pE��-��襖}Y=��"����Y'sq��k`��>3���Բt�Ɂfqb��#$Y�IK��͚����fCKR,�(�<s�5��s1x�;Ҏs�]�=�Nd��Jm�D��Q����˽/t?���(P��K'�a%���^���ǒ^S��),Mx1�����qm�)�^i|\�ֶ��<F�,�	��8P��,[9�8
v50�f͙ޣ�L|��'#}$�)�ԟA�$���2y���R:&��,oe%ԑ��;�j��\�EiR�[��͊�5�F	ݙ�a��)�3.�k.��Yb���,�2��/�X�J�Ժ���-hV-i�Ƈk��\�I��E����S�ޛ���[����kI��,�9i���s7�$�`��iS�:$zK癭�M'�*����yt��?cz}��-�G��8��xڋ��a�\�RS��������(�Wɭ�F��$Ӊ��Ǌd`��4��hL���6L�V�����%�r\�nhd晙�y��>��pf�d�*Cw��\�C�O,�yK��d�	�Ʀckqh/:�k�4�pK�Fgҝ;�ZIڢ��-����ܑN$���