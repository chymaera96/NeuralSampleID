BZh91AY&SYђ� 9߀Py���������`� ^�    � �`�2���ʟ��&  �   `�1 �&	�!��L����  @     �0L@0	�h�h`b`�!44A4ɡ�&��G��6�~$+�"Ze"4����h�	K{�O��
�UJI�E�'�U~�K��">ZFjA��Rz:xW%[�y|�D�b�榏3,[��֦Q�g����G�OWt��Y3f����+:�3��I�<|j�����Y��s9����M�+��౑�;��z͇)|�lV*�V��w(�˪�T�Q8��Zܐ�O"h�����j�Y&�)B����.���لS�X{(w��Eٰ����]mo�Ng�U���3S�%ԙ*���-��
k�ׄqRq�w���ncm��fe|I�X�pSV[�=6�9��0����ֳ���[�_M�����66c</M�n�Y��^����~ř�S+p���ۆ��N4�\n"2B�S&�)b �Rčr}�qk�Y4�e7p�V�4o�p��m��L��@�!"   0cI�Yck�l�#�
>
F�>Cֲ�]E���]��ԣ���m7ԕR�m{UZ֪���V*��Kc5�hɣ%�r���7*E)����ܻ6KA�Cu'��آ�o�ݹ{���������Ӟ�������?�SW���m����Iw��}o���Ѫn5T�M�d��]U~}�ر��Շ���{0��O�:���Jz��|,>�z�j<ʑ�Š��F�ƧΝ���0{"�����?�|�u�^W�Qs�H�$d�����R��)����9���i���g_��Y��},)"��,�Fy��9UY(�z���;>&�
;�d�ŝ�.2T�g��%0޳F�afU���7"�)G��	�A���d��IGa�0��T��6�R�d�f�d.~���C�~N�B�h�����C'��v�LJs.�K}�Ds|���1ڞSg��v��ǁ�6�f���9�K*�Ŵ������~���;��ZL���f�k�G��=�J;�s7�I�R���7=Ic��5laILCМV���jR���)N��j�N
��J.��N��{�♣CM���,RO�w���F��h�cʕ%��ZQ��ji#%�^g��"�s${1�?�����I�#���I�>�'��>�c��vE�:��u��u'D�]���O��T�����/#Y�Pt{GIF$`�_�Ԟ�G{�q�7�ho�(¨��T�*J]aejs\���Qۗ����F��D�#���jf]r��wcY��I�83d��g[��Ie<���u����j���Nmfo�R�
qv*ED����ό���,��FL��D�;Z����&T�sLgF����=-$�(�#gh���H�
2B� 