BZh91AY&SY�Ӄ� P߀Py���������`�T    s F	�0M`�L%4 �B�(4�@h4  @ s F	�0M`�L5?U@h  4     �& �4d40	�10T�hM����i�4hd�2m���I���$KI$�$g#��5���Kx,��E����YR~�*���a�R#�H�D1��:N���ܫ~O5�`7�M8�p��tI"�r�l`Gc���D�\�װ�2�%}��A��Jq�ܳ,�2�uX�kf�����X�߿��4c7�R��zʬ�%�t�e�MK=d�a��"64�K�cZv��w�۵��Y&���UU���yJx(�w��$�j*�ao��,8����^8G�0KwK�0�!����Q��mhԌAX8m;%�Z�bͰZ��Pm0.�&6gY5�)ʎ�|�mcy(;l�_�Śr�A�U'�B"��#���W9ď-*���7q1��K$A\X�!��L�g��5=몒�T@e��
HADB%]��4�=����J]`�E���G$�H��N���׍P~�5&ZS�!B�   L�Z{"w?�G�.Y֣�MjzJR�Qg�c���Z뮲�J���Y�}�H��&Jőb`�!d8�Ι�eWt��(�R�Mj�Jk���k`͊�bP]��d �"���x���ͦ��.�O������?/w�����Xޘ9���?ړY�R��Y��b��U����B�F��އ'��'�7���t�}�����jED�"�X�#c�S�N���>ȧX~���dJs���B��#퉋ě�>�*R�E1t�GY<,j���eU,��d�.��+rge���U��60X���b�5��J.�b�L$[�������%.س6k.����gqG��1<bl3`���]��GA�.�O|��4�6ɪd���`}�޷����(T�7,��	.�8�b���y%�82��ك�����lqN��G���VŶGY�iœ�'2p�%�Ib����S���;6l�j�]Q�ZL����N.��Q�Q��<�N�),�[Ж7����ԑ��;�j�K�pR�Y�����c2�$���tA��2�#2�F��]e�(?����C)��5��-K��=����F�b�g�O#�j��\(�c�^O�%<��Nf$�>�{`����gD`����S��9';'cE='J��Ya��#65H�X����9D�^%Ϲ�������k=���6��]TS�;'b��,,�G�N��Gz�M�lkbM1:ؘ�L�����dnoM���T�V�������K����s���$�0|Z�D���d�U!��M��H�'�T�}EΈ�ֲG��s5��m`�-E�[�a�R8%�3�IN���yT��������)����