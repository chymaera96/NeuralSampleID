BZh91AY&SYSV�3 �_�Py���������`     s F	�0M`�L5S�)�G�@4     ��b�LFCC �#��b�LFCC �#��b�LFCC �#I!0�G�dj`	�4z�OI�ъi��0�]q"�1�g#��E�`%-�Y?������ʓ�^����I��G����1��:Nܫ~n�qtƼ9S7k�-��֦qY�w��ͭO&̴TƱR����[�§:����+��-W2��t���U�MۮS��4�͊�c~�2��̓Ά�tX!��;�cD�&�����r�V)��
����wi�O��LM�oUC��9�e�+�e蛝LY�[��j�,��K+S䴍:�&ʎ���6�Y�z�Y�L�sdPؤ��S�X,���S��˱]�[��g����^����X,,Ä2�AFq����@�Q�HI��ئ+j���e��޲z]��)JUmUUUUUURT���;�7�0,�Q�T�)�<�YR�,�,`��l`������J����^��a{UH�I��-3e����֩��0���ٱZJ�6��u*R�����w�����~�3��������1=����V�h��,oK��)�~<_\�&�EJbԳZ�*���ڋ;�0z�޷�Cq��n�ƞO�>��<���T�"�X�#c�Sҝ-��0=QNH�������آ�T���_bnT����0E1w�#�,�Ve�5(�,��楖|�=��Ec�L�,�sq��l]b��N�/Z�hﱱK�Y��b�E�1���fL�.�fř���gaG�ᘟi����^�����:�$���)M�i2{�b.~γ����np*3r���/&��/l���0��]��&˱������c�vMO��x[�G��ɓ�8��E�Ib����S��~ٳ=j9��ⴙ9��D�NN����%���Rv)H�2Mo"X��5)#i�;�jтW)QF������Z�3�Bl���v�Ix>O�L���Ca��,��'�Z;�2��0�٬v%Ij`�.�3KB�4V-�+;_{H���s����O�%<M�'B�I�=��k`���gL]#��WYN��8.��jS�w�$y�獱�4�<1U7�s��&�����3w�g��9��mF
���S�u�)u����r���.��=_ƥؓV'SI�u�SV���#sznN���ZS�sqIe��8L��6������qf�d��!���J�T	�Kϸ���H�1b�kgWG&��ְ�bƔ�)�Tf|��)ܲ�N�$jt1�]��BAMZ��