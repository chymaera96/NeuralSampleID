BZh91AY&SYR�  ߀Py���������`� t���@   `�1 �&	�!��L���觑��P �     ��=Q��       j~�F��M  !��M0&�у�0L@0	�h�h`b`�"2M�����jh��'�7�6avHKHLa�����	K}O��D��/
,�?5���^!��G�������w�������"�y2�n�,[��-L(ⳝ��5�����&
X�������N|����س.W2��X�ll`��M���\�,�L�|ةP�f`ᖌٽBn�� �SV�$7F�񦋟o�۵T�(R�UWc滸�S�F���{-g*KYX:�f��DԝIL0�r����=���vY��&*YZ��ẛjM7Zj�ڦ7jyS~y+^�Z2��2�=2T���Trt(\�@�U�A)=�/_T'��D�]IkqK0��^q�F�='��H@M�����ka��c�	���I��dB�J   $��^b]�ѣ�sQ࡭OA��.�Ϛ�@�T� �� yZ�vgv�J��Ӻ���.Rh[_KeMe�.�֩��1�[Z�ح%t���G:U(p�q�Q#y�8䭧�m��ڸ�p1\︙ɊZ�~�ڵ�G2��k;�>����f�5�*S���;誯���j,t�h��u�ov���G���O?�O�y�C�Acҍ��O�:[�`{"��a�,�!N�'k�(��H�!����?g%)LLE�T��O�8jQ/�Q�zie�&O���(�qɜe�;��X��b����,^V���'Z�L%�NeF*�,������3f�v0v��\�֋;J>�$�����f�:�g.	GI�0mOt��5rR���d���\���S�����*FnRY=��a����9u��K����v1__��ɺ9'i���S�ض��x�\�:�ŵ8ԋ*�ų����kZ�ٳ=�:�Q��'Y d�'8{�'�IGS�d�);T�u2Mo:X��5)#q�;�r�0J�*(�uR��q�XŵRI�J.��%���%2Ff�
`��O��x�He#\a�X�J����]�f���h�Z��ϱ�Eu�p�=fuI)�pM�m_b�<���l���{�t��:�4��t8'Zt.�v5)�:�$z�����$O$UA����p0����	�3x�Z�[dr�܌E/�d�RR�+C��'8��X��65(��Ě�9�1�\�5k�i��	�6�b����oo),�����͓�ff�f������qf�d�!��MΕH��}R��0:cF��8�-�l�n]�NnŇ�4�qL2�3�N���-$�QRF��f���H�
 �C0�