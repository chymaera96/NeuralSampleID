BZh91AY&SY�2	� �_�Py���������`� �    c�0L@0	�h�h`bc�0L@0	�h�h`bb)�'�� 4���hh  9�#� �&���0F&9�#� �&���0F&
�@#D�� M �P�G���i7`+�	`��G�?U�����d��0��T�qE�'�U�%�f��f�$��)<����V�^/&��e^<������E��sY�w����OF�F�5詚�(��V��9S
f�wuR��ExVg��s3�m����K��n���Í�2o�W�q���kgQ�����FǮH���Hl�5�!�6'�5\����M��j)B�������|�la询��~��xd�����׺않���9-�4�a^��`aIuY_�.gPm���*eR�b��Ujy�v,7)�M�)�f��e���Yu˪�`ݳ�z)�Z5ZR�q�ʭyY6�J�0���#]���^kbV{�V�|[f� ��� �*�Fʥ�"$d�X�F
&	y]f�����w���)U�UUUUUUIB�O`�~m��gj���e=%)R�,�V��u�Xa��ZQ�d��R�>V�cL�U�Z�/����jVK�ͮS����mT�Sm�kj�-E��rxi*��u&ݫ��W���?ݮ���zda���C'�����_5�6�W7ic�]���c�s|�j�MU)�b̘;�誯��k�:y5a�v=/n�a��M�Ξ�y>vt=�x�?(�=H��)�N���>��R,?B��S���~�;d��d������R��)����9���V�آXt����K,����Ee�m#<Ǖ��U��7.�x{�K'��d�1b��b��;WL��w��%0ܳ6�af�366����2>cqh4U����Q�z7��$�M�JS����j�����a�}p�>]�#GT�OIy0�8�}q�S��1)̻9,M�e���u8GRw���4�-�;O	����soNt�*�Ŵ����{j�4=�;<�-&nÕ5:�����%o�Τ�R���6�	c�8j�aICʜF��J�,إ)��ܱ�ި�t�]<��%���%3F���)��X��h�3��F��h�c�*KS%�Ɖh]F�ɩ��cW������c�}a�?����9'��]'��_[p��+�Y�H�<��)�䝉л��ا��T��,<�;r4\k"x�ǸvF�����h�7�������U�J�ӹIK�,�Nk�x�uYv��nmdM�����2떦ͽ-Fg$��l��Y���RYGc��Vn�����q]��\��'6�7ҩ?58:U"��'�^y�1�j��L��Z#���jbv���L�H�΍�:�yVZI�QRF��h�]��BB��'