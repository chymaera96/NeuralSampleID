BZh91AY&SY���G �߀Py���������`�@\��    s F	�0M`�L4FBjz��4M4hb2i��d�&M0`��`ѐ��&��T�J��Sjh �      ��b�LFCC �#I@�h��i�SF�I�ѧ�i�I�b
퐖��B4����i	Kx,��F��H�(�����1j�B��"=t����ғ�wU�;{��t�_���ae�~�5��s����h��t��/E�+� �MR��	�(%�~���Q]�9k���ת�1uۗ]��Uc#vw,��Ա}�S=z���1]LlTϟ6z���A1���Rw&��w�խ��f��JU^G��v)�Y���]O��b�����}g�jT�����h�MO���V�o��d� ��Z�Q�S:b���[��+Z���^ʾ�zs/{̍�-�c���1faL&`�Ф�J+1�P��X�W�Ϡ0 $&�(x17K�	��RD58=�#4�`aE����$C$䔐�H,���ط0%�g
""."����dD�a����e;c�M������(0�V��la��.���R�᭓�%��C)�5l�)8(XY2�H���HR̬�lT�SeSZ�-
��TU�� `ȩF!���6�n�)��e?�;'������+�즧ac�]���k�qxhԛJ�ɭfL�s�W��k��:850�:�������SΞ���6t=5*��Š��F�ҧԝ��0}qNH�����;���\�>�d�&�O��JS�BΚH�'�AmkT�J��q���e�6os
H���6��p�o�Ed�ͫ�^�t2}�'S)�X����݋d��<�f))�ՙ�X�0�Y����wx<�#�KI4T����r��t���s��JS�MS7�FB���0����?�qB�h�%��^L#�;�=��S�ZbS�vrX�n�#���0��I�bk}�)�m[lvC_&n�qnN5"ʤ�m'��)�ؿ;F�j����V�7Y f�'d>��$���3yԝ�R:Y�ǡ,pgMf��b�̴�%qR����j)��ڱ�ܤ�l�];�:��|�f�5L)��X������r6F#F��RZ�a.�4KB�5+&�Hd���}�Q��u��{I�*IO��7��}���>����}泽�Y�H�<��)���iλ��֧��T��,;�v�h�5H�h����p�b>��pOGSsa�m�A�b9��QKĩ�;T�����q\���Q�.ϋkZ�����#���$̺婯gCT37�&��3ek-T�oo),���ɽ���hh�v�����qh�}����3�R*G�L��L��d�0ɓscIˣ�Q���Xxdʔ�)����S��z�I<�*H��M�]��BC��	