BZh91AY&SYo��� U_�Py���������`	? <sZIJY    ��b�LFCC �#4	�SP� �  �  0`��`ѐ��&��OB�Tڒ �dѣ@4dѠ2��s F	�0M`�L$!he6��z	�ѣM=LOI�m&�$EvBId)$M$~g갑�J[��TJ�R]$(����b�V��5H�E|�*!3��U'�����>,�.�����6X��r��
:u]���]M��$�
X�����K)�S�*R�;��Y�]��f��l,�r�l�X�ݝ�.Y�����{&C��*l���DI��{�I-��ѩ<)�s��5kied�$�(UUWc�Y�9)�Q����\_^�ɖ�bVv���� �V`�H�j`�әnWL������詖��CgP��N���Jfq0�Q�K&�S4��)�V,�Ă3+���9��U4fdC���PmN�TOxjF�Sl%��@�4HQe.��M�5�Su�݄�f[���5LS;Ő�V�s4�l�a@؍7�X��j�"��u�T�)���H���E����J;va¼-a�cP��<�P��oX�ϖ�x��u��	(�*��L��4j�٨֎W-#����9��#5P�j�܈��9woA��{k�3ʂ�B-�����Xԋ-$�4���X6��@`_@��b����)�t3�y��s��J�'.:W����&�CKIõ��:�kP�n�j{�Sm[�Z�qb50�w�i�C�ʫ}�v	e��,e�E��-oL�E��N���Z�K�0�UV�7�� �00�s4-t��S��E�E��Yҙ�������]�B��  �fbU�=)!����<`��j��SaO9Jii�J0�V�.�c4�u.1�T�&!�����Ή�$�1[�I�%E�035�v��I�P�A$b��c�x�i�.����"��G��ֻ6KA���O�7�q��@R��Sf����no�׬����l�t9��Ú��C'������E��SS���Ηnix���p|�jM��Jdֳ&�:*�����<�L=OS���H|#�����'��퇘#P�)$?H�;ѵ�Sԝ-��0}qN2,>E��jHS�����.u�bHd�z���)�S!g��8H�|�5�,�T��g��Ygɛ�(��ͤg�Hw7��Y(�j���:Y>�œ��K�h�,�YBL�	g�
Ja�f�.��;V����giG��D��ZI���'��Ε'��r{d�	����T��Q����=l>��{�P��d�y�ɄyGs'�?d��1)��9,M�e���0��)�bk}�	�m[lu�_oHm��AU%�i?�N���4hz�rꏂ�f�s�Bf�ZH{��\���f�;T�x���K�ᩬ9�C�9��W*��,֥)�q�X�nT�m���v���Ħh��n��)��X�#�-L�3&��h�c�*KS%ޖ�h]F�d�h�,jx�cTEr�9$������T��S�7�F�����{�������gL]#��YN�:rN�ܝ�jy���Aa��E�CT�㊨9=c�Hs�Ik�9��h�nl=-��6�G20��^%N�ؤ��V���N���,���j6�2&���F\S2�ũ�gKRHfos���f��Z�����QɃý���yu�f������ph�3}����S�ҩ���^y1��d�	!�&�Ɓˣ�Q���X|�eJG�th|i�)ܲ�O��5�G�rE8P�o���