BZh91AY&SYt�  ?_�Py���������`�E�J�   �0L@0	�h�h`ba�l��xQ��      `�1 �&	�!��L����@�        �0L@0	�h�h`b`�!C M�Ɂ'���6�'���6�v��bI�#I��,��)o����aQ*�RH�(���ת��Iq�Dz)�A��Rxv��*ߋ�ɢK�+:h�ſ��ja�Vv���ty����m�M�T$4�U]�bV%y��T�q��o�]W3��wX�ons.�3z�G�SY�F���vX�e��{gV�S58sٵ��"sC;H�ѝerC�0�$�q��v�}k"�B *��xe	�!iI
tW��w],�Fr��T���]��{�4��k��+�����7,��Qz۳E�ṋ�}�kmY�K2�K����J��ϱc{]��*��5q�Z�7�u*͙�Xa�ٮ�\lR�$��% ��k���$<�L4�d`B���$$�dDӪ��$�扪���m����I��L��I|�ң|Ѷ�Sc���v�IM�����m��nk㵜���;�JR��UUUHB$���=K�h)	2�?Tڧ�R���?E�z]��YE�'�F7)�eER�m4^�c�^V���(`Qa�efeH((�.��)�Sb�Y-Ei9���U�u&փ0��F�?���F ��BFG����m5qv�9���/���T�j�L�d�ܧEU|}��ac���S��y������<�q>vl<�55�Ac΍ϥORt�?4��rE�ĳ�n%:��آ�l���'̜?g%)L"�:�#�,�&Ś�$�J��q�y�e�o�(��ͤg�<z��Y�u���N�O��d�Q�p�k+��ݫFJ�0�A����f�b�,ýfb���Y�Q�y&G̛�BΆO˝(�<���$�M���4�������������8:
I���O���G�x2{c�N]��N%��bn�(�/WY�'4rN�c�qO#rۣ��93u�zq��U%�i?wN���4h{vuǽi3v�C59;I���%O!�ʤ�R���6��c��5l0��c�Ne�a)Ĥ�͊U+��ر�z�n�����Ix>�Lѡ���
ae�*I�-l�3��14X�J���	w��ZQ��jhL�5x�[X���;	�zLI��IO�Μ$���]'������gL]#���+��C�;�wc��O��T��,<V�h�5�<�Uc�;	�`�>��s������z[��n�daTR�*wN�%.���8�Y�틨�o���F��Dّ��˒f]r�ٷ��389ӂof�VKS���������CE$�.�5\��'�7֩59�*�I?��e��`�[VH�L�7��I̺951;]��&T�qLgF�E<ZI�QRF��h���H�
�Q$ 