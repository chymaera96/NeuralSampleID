BZh91AY&SY	p�e -_�Py���������`�xAO^�   �& �4d40	�10��?Jm=(  �     TƊ{J        	5"����=i���  �@�& �4d40	�10T� �h���LM54h1&ji��pB�ȖH��3����b0���O؅�Q���!C'Բ��%�!$� h���'_�c�5�[�,Mn͉�ar�
���.!�(߱����LmCu�Tˉ`A#���m����	�NS�����s)��e���m��7UX��h��ڸ4��`φ�zRٺږ_�G�	��!V�rC|h�D�s��{w8�VI�)B����.�|Tj����xvcM�^�b�S/\�ò�9Z��&�����P�� �C19��u\��z�IV�%�����{冏�1�*21��În��z��/F.k�ig.ֳ�i����0�i�A�A����nyZX�&�

a�C:^�	y�ϻvŭ�5���2�lY\��p�ైհ��|f���8B��	аa`�Z�7-����8�b����*���HQS�CY�i6��GTC�&q6�#(B��RE��.\�
�fl�����I����DrI�.^�4���PSQ�R)M�c>���1ZJ�o�E�I�e�x^Z��9t3���.f�L_ǋG���K��M�Ŏ)v�w�}o���D�h�LZ�Łާ*���]�c��Fk��{�np��G�cО���+��h<�G��ǩ^u>��m~I��tE��Y�����Ԣ�t��F/�8*~��R�"��:�#�,�q�C��}~�Yg���0RE�93��G��ƫm]b��S���lY;X�P�ڼ�qd�Iy �RSՙ�X��<d.j؋<
>/4��#ih3U����N)GQ�0nO|��k�Jo�I��s�w�>�����P�f�%��/&�/|��ژJs.�Km��s}=����<&���<ͫm���kѓ�ۓ�ʤ�l���)�ؿ&lٞ�����'iƐd�Gr>��$���2z�
R:�&ǥ,qe�)#y�<Sz��+�����T�8�{V1��$�d����^�����46�)��,TO�h�e!����f�c�*KS	w��ZQ��hf�V4y^���v����I�U$���"7/�t�#�p{�G�jx�:����s]e98�jr]��j��u�H�����$O4UA����q0F���)�3v76���F�*�^%N�ޤ��V�5�;�u1��Z���Ě�w11�\�5���S�n�1Z��N%�v�<�2r���������sf�{�!���R�Q?t���9��6,���nlfM룣C	��X~���#�a���:�x���ʢ��[�����"�(H�I2�