BZh91AY&SY��+� �_�Py���������`_      `�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L�����`#@�#@ڍ6�4M�ق+��d�����0��,��F
�UJ�]E�'�U~�K��*Dz)*,3�������a�t4���e�~�5��Vu]��skS��ў>k2S�J��e9���S���ՙes)���ca��r붛V18p�f�[�^ږ]{x8kŚ�D��� �իV��֝��s��n���Y&�P���~����>�50sг��wX�ũȷ�0T��9��SQ�?cT�Ie&R�W�LJ�F�f��׎���%6���0s�SR�&+'j�so�i���o�n|o�eζ*��%���&&7�Բ��*�ک4dͅ-�����i[�Uk`�wu���U)JR�b��������Zz]�ћ�t����O1JR�,�V=�����X���h�,e�f�᭒��*�R����kUI0/Q�R)Mta=MK�1ZJRn}�Х(�I�Z�{kw�k���>:�\��|`�O����84~>ߪ�Z飋���.���O{�q}3h��)�R�XjsUW��k�9�4`�^�����n��<�y>�l<���O�-�:6<jz������)�2��Ng'k�(��$}�_RoT�ܔ�0E1x)#�,�E5+J�*9�G��K,��{X)"����Y;��X��b�����^&���F�-�WS�.�ILd�b�`�Y����v�}��l3]9��\�s�`ڞ�'2j�7I���Q�����������(��K'���#�;ؽ��'.��S�vRX�.�#���`�����j}�)�l[du��L���E�Ib����S��~flٞ�=�ZL�'
D�NN���{$�x'�Iڥ#��5��c�(h�`����M�%qR�Y�JS�Ǳc�	�J.�����?"�#3��0Ye���h�e!��q�f�c�*KS	w��ZQ��hf�cGs�i]<GK���I�$���7�ھ��}O{{��>�Q��,狤t�I�u��pN��]��jS�x$z�����D��T/`�p0`}����C7CkY�l�A�a�����T�jJ]aehq\���Q���cR��lI����$Ⱥ婫_;FF�ޛY*����oo),���ٽ�'4��G��w���(�Y��>�Ho���Ω)㗞3�4kY#�-�l�ˣ�C	��X~���#�a��*x
w����EI�I����"�(HlyԀ