BZh91AY&SYG2]p ~߀Py���������`_ >G�5R�(�0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��T�U@   A�   �B*~���z�D=C�='��@�h�=@T���jzi�����4��4����	+�Y��4�|���K~����1)
�*H�*,��~�b�UUW��$���f��,YP��y�+�ww��uC*���Ybߗ洣
N�i�]��
���_%���cD�E�%_�;FJi(�����9ܮ����Ϳ!��6�c�X����B���I�\��83i/�V�&2ٴ��Xv1�n�v�7���-$Sn���Ms�R�<��(����vVcR�����]�N�?E0�N���`^4�&5H��̆�L4����:w���`�P�a�O��$yn���n�H+��n��i��+9˕d�:��d�jj�aˡz�cE�Z2�ŝm�̙��k�v�Չǎj����%[u�錘V]�Y|^VLm:����9U�o]C@�����L0�T�!H"� UUB�->c�~M)1T�c��7EQ򬱭����JZ2|��^na��*/3��U+�m)u"������/F�,���s��̭{�_9W�^M�Jn�盥�̖D�R4����U(��Pݹyw�\>�_\�f�s���8O�L7Q�zJ�M�W��7���^�ˎ����qu���6�*g7��GqS���?��m:��9���q�7���Z��p���6��(��d���ޥ/쓛y�,a	�?���9��^T\�[�[�8@�0@T�5�#D ��?V�TF�VR���:���|�X��3}L*$�Ye�I3���N�T�M����KE�}���7��hw1h���g�~���*$��4RT��Y�B�v%������r,zE��̓��%IgS)ޝ��I�<�:!��қu�N�g>�J�;`���R7�ݫ)��. ���PM
k�Vy���m+FD�ZY��I'[��`�8GX�M�j��'�o��'q�u�;gD�u%���~�h�蛗�4hi�I���Z�S�H3)�|G���(��g>B��QQ;�$�rfMM����28,0��JJ6.�*���=�I�tJ�^:'R]#�{�gA���L(���qi<�4L�t��F��|�/{/%�<�����j42,j�:cFh�Т���Hu�R�v����[����'��:�����ZS��;dt�;]͔�;
�,��ˢ&��UH����I㑑�g�`����ZB�Ρh�[�)PD$*y��R�Y['Z�gk�.Tve����J��RM�̓.�g]-F۹�����#���͕-ij:�.)D���`��53:f�hT�#�w��s�C�����)��Q��T�����^z��MM��9��6g�����F#��Y�R�֘ΓI=�<�O����h���H�
�K� 