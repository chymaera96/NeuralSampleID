BZh91AY&SYU� �߀Py���������` �    9�#� �&���0F&9�#� �&���0F&9�#� �&���0F&���        `�1 �&	�!��L������4�@ �#A����4�M��RE�bC9����)o����`��T�!r�*O�z���K�%H�E#%H��a�'�uR��v�d�N���L�,[�|��qY�w��f��2��R��y0��<�v��)��+���+�L��,n6.�u�[)V1/i3n�nuJ��b��M/����Hn��HCkLv`Hn�I�MK���n���̥
����w���F�8�����u:�/ѕYx�s3���,�*�*��g�x)�Tg�e�5�SZ5�)j3UՋ�j�ٌ�F�-���ě��he��]ӥ]KZ7���db�YT��Lhk��Xn���*d`�{,��n̚��mɌ�J�מX餭�jTa�Xe�wa=F�!B(   Li4�)6����sQ�Q�S�y첢�,��`��l`��J[�;�e��f[*�*��֕{Z�ֵPfŅF�H�5ь�5.��h1(j�������(�I�Z�{��k���>:�=϶0k���b�\?/o�v�t���X��mgx����}3h��)�R�X�tUW��k�:x4`����v���n��<�̟[�T�xT~�h,yѱ�Sԝ-��0=qNH���:��آ�d��1}I�S�rR���Y�IQd�5-4�Q*:YG�祖|�=��Ec�L�,���V*,غ���'K��f*:��\��;
�Ix �RSř�X��;�d.jkE��G�1>���5"Ά/˂Q�yLS�$�M\���4�>
1?gi������;��&nRY<���A��������K����v1^��&���S�qO��m��x\�:�-�ƒʤ�l���)�ֿC6l�b�}q�ZL��I������{$�u>�'�Iܥ#��kyR�PѨ�I�!ޛ�L��J�5]T�8\{1�U	�J.��%��ߙL���Ca��,��I���RH�Fl�;���0`�zY��u+�f+</kH���s=oI���RJx�|�j�I�>����~���Y�H�y'�S��9�B�n֥<�R��Aa��6#5�$O�*���g�~�����Z�Kdr�܌E/�l�RR�+C��nȺ�X�|[�lkbMX��Ly&E�-MZ�Z�zm�*�����%�s`x7�d虙�<��0D���d��C�MΕH���/<fLhֲG-�l�r����v;V<Xґ�0ʌ�ҝE;�ZI�QRF��f���H�

��@�