BZh91AY&SY��W �߀Py���������`�      �& �4d40	�11�& �4d40	�11�& �4d40	�11�& �4d40	�11�& �4d40	�10T���&�50�L�4P��M�jj{Rp�+�I!�CB��i&!)����T����E���U���3T�=���I��Ry��j�W������/'�^m*m3aih���,��v,��?-R�Y���b����,�Ч}U+���-SM0e3;{m���q8����,�����]��;Y���U3{"8Å�Hn�m��7�G�M������N���MJT*��ߪ��O���%:�v��vVt��4���4i,�Y�;���&��df{�ڦ|"J��k-��8�ڝ�NL2�i���#3vܳ�LT���u.�gB̩9JR��k���ݫ�v�6r���YQ�:�[�e���[�F��-,�m9f͆U��ݍU�j��w,���j��u�xy}�R��*�*�UUUUT�Yi�<�G�1w�>�n���J��~���]v�0���e}���u��++Z�T���UEYhY�̴,�Y�UF�%)�F'�U��Y-E�NO�;�T�*M��]�+�����k�=��NO�0ޟ㩓��Z�/��m��񖎔��4�S�?�7�F�%�S&�2`�S���O��شu��a�w=ϳ.���Kw�zd���>��⏭5
>Id,z�pz�\��&rS��g�p)��W�<b}�O�:��픩L�L�g���E��ڤZ٧��K,�ϺaRE�Y�#<�C��d�
]e�/�9�y���wJ�3,[��-2P�y`�T�Ä�͢��Y���1sf����<�#�p�!��:�<�gJQ�z�8��I�b��5��FB���1=��G���ߥ�)��E������D�|�����싳'�H����$�Og�s����,m���sqNt�U%�i?w1O��4�4��Gw�<���I3T�x���{�}FoJ��JGl�7}ih�f�[P��#�'%�	Nr�QQf�R�7��c'p������.����F��)��Z*O���fFr7LF��(�ja�w��Z�j���,j�l�"��������AO3�:$�W�O���s�?�ly��iq;��9ˬ�S�;��ws�����B{;���#V�>��C���Q���Τ��;�[���;d8'R2U�J��IK�+c��i�4��̼�����D�#�22�L�˖���jft:�蓋9Y,�Y��t�Q����j��44Rz]σU��sh�f�TGG�NN�H���藞�Zj�a9��6nS�T�'kh��y�L�R;$�th|��)�Y`��P�N14���)�8�B�