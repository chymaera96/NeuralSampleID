BZh91AY&SY��c� �_�Py���������`>|���`    ��b�LFCC �#OD�Dh� 4  �� �  4      �?�D        "�(a��4i�F�@hd�2�T���� �� �SF�4�=��INu�Ed��J����Ip%�Hs���D(̡"�"?�df��f�FVXiI���[�o������e^<������E��qY�w���u6yt��aKRQԲ����S��Wr�Z\�fl�cq����dnX���fL4y�yϿVjT�SSVY�ѣЃ��l�5�!����{�72�XL�)B�������|�j�)��=x�p�ÒT�ш�@Ba9,���SS56�Vl2f�)�w���uzg��ؾ[����x,��3R��|�ce7U���P�[��#�;���MZm�����U�L��F��WY�˫K_9%�U�Z�8Xc(��X,4�4,EfLA�3e��fK5��1)�ֺ�6k���j�#w���T��	H���h�EeI�R�j̼X�*r7Y�	�
`�PiB�f��ha6'�2ʠ���ť=� �� 
���-=2���F;T}ڧ��)e~�Dz]��YE�K5�jJ�ZZ�V���|鱕�J�Y�ey�K*�^�Ihک��3���ٲZ�i9��C���(�I�j�{k�k���N;}]w�0�O�����5~>ߢ�i�����.�ix���q|�j�MU)�b̘;�誯��k�:x5a�v=�>��|c�k��O/�O���,F�ĩ�-�:7>�=I�����)��g��!N�'��\�>��BoT����0�d,ꤎ(�|�Dl^,��祖~���Ee�m#<�;��Y(�r���:Y>�Փ�F�X��*'j�JH��B��nY�E���
��͍���Q�x�G�Cqh4U������s'�IЛ9)Ny5��
2?gq�����7�
���K'���G�w�{���.�ħ��7]�G��Ó�9'�����S�ܶ��<�L�R\�Ƣ,�K�~�"���4h{vu��ZL݇
����!���%O�Ȥ�H�f�^T���5l0��s�Nu�0��JTQf�)NŌ�ʄn���~�Ix>O�Lѡ���
ae�)#�-l�3��14X�Ija����-��Y54��cW��5���#�C�����T��S�oI9�ܺO��o{���l;��1t���8���	؝�͊y��I�ý�nF��k"x�ǰvHp1!��~���:�ͧ��9��FE/�t�RR�+S��nغ�Yv�[�nmdM����&e�-M�zZ�fopM��͒�U���%�v0x7�f�*#�޻��s8�Z<L�b�7��t�ED	��Ϭ������C&Nf֑룓S�ܰ�reJG�th|��S�e��%$lsG�rE8P���c�