BZh91AY&SY���� }_�Py���������`��)U
   ��b�LFCC �#��b�LFCC �#��b�LFCC �#	M
i f���� 2 ��b�LFCC �#I �&��cD��SG��#z��I�J�%�C&r?�ZD�J[�d��0TJ�Q�QeI�?D��V��FJ��FJ���w�좾n�왂�QR��8?78�DÝ(9~v!N����`��))��OR��R���W5�p���ե�e�l]v���Lvܥ�<��s��(:�eM{��`��YFl1Ձ!�'�5.}��MJ�X�pR�UWk�]�9)�S��Z���{*J��Ԅ'I4���f�X�(��b�EJf�&YZ˕��4s����{+i�6D�HkFDr�.`EH׉s��h1���j#&��0d�F��#,^�"^MզhT���!3e�Z��9i��y��e��ue�������J�iFQ��m,�!���=k���ʣ�E�D<��u"��L��T���K]�`~������B�%��I	$�0;w��1�����JkS�xYf�e�c洂�d�mBg���a�Y݇N���CܡF�RI���C	�!;�����"��G��k]�����'��f��&�H��k�<^�������bL���b�;�>g��Z飃�cz]���k��xظ���C�$8o$���f�r^�'��kr|okv=)����CA�T�Z��T�����&�)����l��..��Qs�����ț�?W)LLE�t��OcR��I&�¬rwP��N2D3)R�e����TY�u���:������F��d�T9�Iy��RSř3X��;�d.jkE��/D��ai&j�t�y�;Ҏ��`ڟ	'Jj�:$�d���\�]�c���w:E
���K'���#�;ؾ�'I��줱6]�G��`��)�a5>N	�l[ds<Ʈ,�ppmN!eRX�s�p�k_��6g�G.���&NF��d�8>>�IG[�d��;��u�MoRX��5)#���д�	\��(�uR��q�XŵRCd�];�:�����#3��0Ye�#�-��2��0�٬w%Ij`�.��KB�4V-��cG�����\(=�i���RJ}鸓j�I�}�σ`����gT]#��YN���+�;Z���j�=��{�،׃I�Pr{�(7�A��?czx��Z�kdq��F
���S�v�)u����r��8��8����lkbMX�ؘ�L��Z���4�#sznM���Yj�KsqIe�m�:ffj���.��\�e�7���T��%:J�R�}2��0:�F��8A�ֶr��C	�ڰ�ō)���i�S�e��u$jm&o�.�p�!S�_@