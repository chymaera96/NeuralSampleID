BZh91AY&SY%�( R_�Py���������`�@�    ��b�LFCC �#��b�LFCC �#	M	����2i�   � ��b�LFCC �#��b�LFCC �#I ��&��`FLSF�4�=&z��I�+�"X�bH�G�?E�0��Y?���$���*O�z��d���G�����a�'��T��]��$��kl����8?��:$� �B�-�#].��u,QIQ/KT����T��Q]�:x��dr���b�]�ر�{I���)kz����fY}����:!��"6�j�C�5'�5.}��n���hJP���~���5<jt�p�+�뵡]
�r�X�p��8]�x��%�d��]3<ϑ���=�m؍�
Z����%�՜0�#R��Đ948�'Lm�`[��\��pת�5���d)�"�譊m
��z	#:�]K�s�ji	/^_I�O�s���)���`�D0] M�$�9h0�(�o�7l,���4�H#C$b�0^�A��q�B��$�����(�Z{	�������G���#��M>ㄐA�I��'L~*,׌��d�a�'wI����@TEIr�:LR�1�3FPCr ��P��I&a5��� ��#ƕ�4ώ���������1=����V�h��,oK���S��8�3h��)�R�X�p����k�:w�`����~��>Q�����'���BM�D���X�#c�S�N���\S�,?2�ᰔ���~�;$�q1x�r���)�)����8����5,:YG��K,�پ�
H���&q�D�n7�b�͋�^|�b��b�:�إ�-;
�b�E�H1�űfL�.�f����gqG��1<I����^C�����6��I�5rR�i2|Tb.~��������(RLܤ�zKɂ<㽋��r�Jq.�Ke��q}]fN���S�qO3b�#���2u�jq��U%�g?wN��3f�����%����D2S���Q�Q��<�N�)L�[Ж7���F
H�0�zt,��*R��WU)M�Ռf�@�%N���|�2�#3��0Ye�������R5��5��-L%��ih]F�š�1X��{�DW>#�>���O�RJ}�Hھ��x�罰}ƣ��Y�H�y��S�zsN��Z���J�=e�{�،�&�'�*����d�`L���������{#�lGB0U�J���IK�,�+�u�"�9c��ljQ���5bv11�\�5k�hL���6̕�Ҝ��K(���nh��ff��v�����qf�{�!��N�J�RO�>�y��1�Z�I�ֶi:G&��ڰ�ō)S���Ө�z�I<�*H��L��]��B@�z,�