BZh91AY&SY[�� �߀Py���������`�<����   s F	�0M`�LEO�E<  � #   0`��`ѐ��&��SBF�z��y5 h ��  s F	�0M`�L$@�bdh�'��ѓMM����OI��oRl�+�	`���G�|�C)o��(�Q*�R"�*O�z��d� ���;�b�ff����m{b~�����*��p��tI"C������f�91�*\������Z��L��S��W�gVw2�k�����u؛17n�f,�Ss�+vmJc�V��4ɛ7�$tCm����.HtF��&��o�۵�eVI��
����w�槂�LNh�8XmƖ��R��L}o�\;ifZ��c�D��,��l��U&�KuZ&N�f;k:���ƥ�56�i�rt�V�az�v�+�A�T4�FiY�6��"�A|(ȭGɇ-G��\�8X��>|n�0]y.��VG$�Â	���D�"Wԅ"i��L��j��7ݰ��$!BY�$�I$�B�OX��oL`Yأ�RkS�z�YK���`��lR�
�Mu����{�P��yx���5�KJj�(Y!�jZ�Z�R���}mk�b��5�i<�T$!Hlq"
���z��V<�f��ĵ����������v�t���Xޗmgx���8�3h��)�R�X�p����k�:w�`�9��^������[Ξ��<l>�z��~qh,z������Kc�L�)��g��)�����.vIыě�?g%)LLE�T��OpԢ^,���R�?FO���(�qɜe��n7�b�͋�^	���5��(�Q��Ź��Tb��<�b))�b̙�]���255����bx����Vpb���'���=�N	����I�ޣs�v�>����s��H��K'���#�;ؽ���.i��줱6]�G��`��I�a5>)�l[dvCW&N�ŵ8�,�K�~�"��k�f͙�QϮ?����@�NN����%O1�Τ�R���5�	c{(h�`���w�B��+����R�)��ر�j�M�Qt���/��)�30hl0S�X��h�e!��q�f�c�*KS	w��ZQ��hf1X��{ZDW>#���	?�����t���.��������5�zΘ�G3�8���Ӛp]��ԧ��T���;b3\i"y��o`�7����������z�#�lGB0U�J���IK�,�+�u�"�9c��ljQ���5bv11�\�5k�h277���Ɋ�U���K(���nh��ff�yۗ{�.`2�ś���T��:*�H�闟I��5���bŵ��:G&��ڰ��Ɣ�)�Tf|��S�e��U$jh��rE8P�[��