BZh91AY&SYЮ�� �_�Py���������`T@	*    9�#� �&���0F&9�#� �&���0F&9�#� �&���0F&�DM5M���� F� � �`�2��*H����4OS2b�=@ڌ�3�M�M�$��`-F2D�G�~�@�J[�d��0TJ�R$��E�'�U~�K�L�"=t���1��:N�\�r����ـ�"�w#'qC?��(�h�RO?�'�G��؈����jً�i���)����Juz��,�빔�׶��kc�$��0� �	Y'P����ǉ4�J��Z_������m���cbBfʱ�!�0N��s����3֬�I"�*����w�槂�SS}}w�I��*�Y-k�N��$Ւ�1*�.�Ӽ��������g���oNd�0"(L^sN��]����>�tmU@����R1"�3/Y�sfnz:!#fe���h�Ef%����04RK6z�	�z�N)0ٻ��Ih�����8������$Dl� �K����֭��g-�4s�iiM���pN)���7U�Ϊ�fb��,R6�ܜN�m���Mp�f5\�r���p^�S̒�k9KW���1w��!B�	$�������-=�Gs�������5��)JYE���z�]��(���38'v�%�K إ�5��ee&1�HJ���Z���	�*ERkT�S]ϩ�vlV�����'�	A�#}ɓ�]~g:���{w�v�
7O������}�g��Z飃�cz]������͢k4T�-K1`v��U_���j,uoh��rzެ[�����cΞ��<l>�z!4UI�Z�l}*}I�����qE��Y�6I�qw?b���t��ě�?g)LLE�t��O���"��eU,��d�)"����YI����TY�u���Φ/��d�Q�$��9���Iy �RSř3X��;�d.jkE��4��6���,^C�����6��IҚ��N�4�>*1?gi�����}۝"�Bf�%��^L��^��S�$�S�vRX�.�#���0qtG�0��'�6-�9�CWN�#�jp�K*�ų����sZ�,ٳ=�9vG�i2r7Ԓ2S������%o1�Τ�R���5�	c{(h�`���w�BИ%pR�Y�JS}ǵc�D��Qt���/��Jd���e�)�Z;He#\a�X�J����]�f���h�Z��h��"+��H���	?�����r��]'��n{���w�+:���<��t��$�]��ԧ��T��,;�v�f����抨9=�����H��_��<ݍ�g��8���t#QKĩ�;T������gc�]Gy���lkbMX�ؘ�L��Z���4�277����Jb�t�7�QɁ��ѓ�ff�O;r�E�Q83yY=ʐ��C�R*�O�^}&ThֲG	#-�l�:G���a�R8&Q��Ӭ�z�I<�*H��L��]��BCB�#�