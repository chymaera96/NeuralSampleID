BZh91AY&SYs��� %_�Py���������`�� R�   �0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`ba)�	F�S��44 4��0L@0	�h�h`b`�!#C M�Dɑ����'��=z���)
�H����5����h�BR�5��(¢UR��yYR~��1j�B�C5H�U*M�;,5����Q_����%��-3f���r-L0��g]��F�+��3��0�
))�W��kݿ&j\�!on�s~�jn�9dT���:@9�ö�#q8�J������l�a�D���DF��ۂC�6'�6��K\�iPk3@$��s�p�XG@��D���^\ii:M�c���%M}o�Z�Sf����~էK[9$��T������E�v����OV"��"�5a��l9��ӣ�I�'N�"2j��Am�2=l�H�9cS�z��vx�HTWxO$�-c�	+�H��Ѫ�Dg���E��Y�F,b����5�LXX�Lt�̞xx2�����n3h��!	h�I	$�3	���ci�0��)ث*m�������)cq���`�"� AFy"UN%�;��Й=&40�!UXtP��"I3�$ꍪ�Jm��bj�c%��CZO�7�lI!3d�"	�>�w�O�jk�L��1#D�y�?������]�m5pv9��F��}����Ѫm5T�M�2`�S���_]����Շ�����r7��ͮ��z>�x�}��D�yU#�Ac�F�O�:��`�E8Ȱ��)���~�;$��FOoT��T�0�d,餎,�6�͋YIT����ie�&o��$QYe�H�9���VJ,ܺ���'C'�ڲu1ֹf��d�v�RE�H2��r�,]��w-366��⏛�2<dn-$�R�y��q�J���aȞ�':l�9d�f���\���������*&�2Y=%��<{'�?T�֘��]��&번����8�c�w�{�y������ś�F�
Nʤ�m'��)�ڿ;F�j����֓7Y�R�����Ol�������R���6�BX�g[)#��;ӕh�J�UQE��W5ǵc)Ƞn���~�Ax>/�Lѡ��S,�I?����C2m�F�;���0�]�h���j���H�cW�������G��1'�T��C�7���]'�������6�zΈ�GY�8.���d�Nu�n��='J��Qa��nF���D�EToh��bF�����4u9O[tq�ʌ*���S�v�)u����rΧd]G]����YfGc#.)�u��ٷ�����dޜ�52������IelM�Y�熦��f���������f��!��NWB�TO�<���`�[VH�#&NF֑9WG�'c�a�ɕ)ѡ�IN���yTT���M�]��BA��K�