BZh91AY&SYbءc �_�Py���������`_      `�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L�����h�I�L�"4��54�Mؑ]�"�2�i#���0%-�Y?�*%U)!yE�'�U�%�5H�M#5"ee����:�U���H�x����l,�o��0K;���u1j�R�]��J���K���T�G���9\�fm��h��]v�c(�b�[c���&Ƭe�R���ǥ����o���؞$�s���s4�d�JP���~��gb�%��s�M��:�I�c.L:�d�W�t�M�b���/w6�"��B�[�T�L�V���o��%4;�]���ЬXl�hⲗYRK�ٳ%�<i{c~yWK'A��gKyvL�յZɖ�6�ƕ4Semk���/���e��*-E7)ux���w���)U��������������<���5M�y�E�R�,�V0��1��X��Z7.m��*�l�E��V��{UIe3[Z�f�I�R)M�bz�h�h2(l���d�(�I�j�{k�k���N;}}�ta���pj�=�5�6�Wic�]���Os�q|�j�MU)�b̘;�誯���l,t�j���y��9���86��d�~�|�>�}1��~qh,z��S֝-��0{"��a�,��:��آ�l��̟2s�~�JR�E2uRGY>M�b/�q��R�>,���Ee�m#<烜�U��7.�x9���mY�j2]bݧj�*H��B��nY�E�������QgyG��L���ZgC'���(�>�d�$�	����&�7�FB���0���|>�B�G),�r�aa���G�N]��N%��bn�(�/_Y�&���&���Crۣ��93uN.d�QeRX���q�m_��F�ԣ��>I���R&jrv�����u>�7�Iޥ#��m})c�8j�aI�C�7�J�*(�uR��q�,d�T&�(�xjt���~%3F���)��X��+G[9�m�F�;Ҥ�0�]�h���j���L�5x�[X���;'��1'�T��G�I̾��|�s��7��x=�:b���q]e:�:v;��J�=%���܍�ȟDUA���d�b`����>F��3i�n�A�b7�
���S�w))u����rηl]G,�~͊76�&̎�F\�2떦ͽ-fg;�s�36V�KY��s��Q����h��44Ty���W03�ţ����C���J�T	嗞SLjڲG�'3kH޺951;]��&T�qLgF��N��-$�#c��?���)��