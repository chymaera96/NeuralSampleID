BZh91AY&SY�Ί� �߀Py���������`      0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��RBe1�dɣDѠ�L�A���n`��I!�$��Y&��'�Q�D��I�YR~K�W��\�D|Ԍ�"ee���N��~/>3K����S'���-���S(泺�㣂��NmTp�e�)+��mz�ʥ��y*���+�fY��fm챼���u���V29r�M�\w�3���f�=����]�Z4Y�Hq��HCsf͘$8���M��O�����Vi�JU^G��w)�Q�a҅�ug�P�TeOV�)u�s���|��T�D��d�����}��ڲ���y^	��k�}1g5��g��vN�a���a��:��9|�[�m���M㍓�fU�+�d�H֑�L�]�������ό��Ҷd�������w���)U�UUUUUUIE������zc��>*6�zOU�T]E���]��0���ѹ�q��־�mXcI����Vv�U�j���U"��F'��v���"����;TR�ԛv�w�\~�_\�v�s���p}Q��~L�ϓW���Wl�M\�ŎIv���}O���T�j�L�d��S���O��l,u�j���{�7����]�B|�i>6d>T�yT~Qh,z���)�N���>x�DX~���qN�G{�(��$}O�8�~ΊR�E2x�#�,�Ŧ��l���R�?Fo��$QYe�H�3���U��7.�xY���mY���]��ab��2RE�H0))��4X�0�Y����w�|i��7.��L�C�$���L7��Iԛ:)Nk3}j2?g���{��}�]B�&��Y=%��=����:v�%9�g%���9���#�w��k�y���ǐ�ћ�soNt�U%�i?w1N����4h{Tv�Gങ�NTI�����=�J<O1�Ф�R��f�_*X���RG�N&��J�6]T�9\{V2��	�J.��e����3F���)��X�?����C9c�E���-L0�z�%�u�&��K����Ev��������IO;�q�o_r�>'���7��x>��qt���9���NIڝK�^6�='�RG�Xx=��sY�Pv����`��?s�|���:���*�^%O�)u����r��t]GL������YfGs#.��u�Sf޶�g$��j�J�S��Ie�N-Y����OC�ﭪ�q9�yY��Hq���֩��|���0uƭ�$s2d���8.��LN�a��ʔ�i������S�e��U$lo&��.�p�!/�8