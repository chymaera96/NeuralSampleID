BZh91AY&SY�[h �_�Py���������`�      �0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`b`�!�C$��4�bh�a�G��MOjM�I^,��!���~���+'�(¢UR�J,�?5��I.�5H�����L��ғ���J������y�?=2y�Yb���Z�aG5��|?-S��шaKRT�ij�JxxU)��+ʳ,�g39���l�ں���\�Sf72���c'kCGV3f�������۷`��'�7.}�V��5JP���~���r��t�g]l���h_��b4�CVw�;���h�%+�:��&�{����t���|���U�ʭ������řh��'������k��s]M�M���ث��Ѷ���M���e3�[r�q�~�ݓ��YSm2��
Y���Lfѿ	�p�z���匪�oU�nɱ}���7�=�R��*�*������),������z���>JM�=g��*]E���]�ae*|t[V�I�V��6fɪ�%T��j�Z�RLר�R)M���6]���dP֓��'}UE(�I�����/���?ݮ���u����j��O����}%۶��n��R]���k��|tj��S&�0x)�U_��k�;:���;���R~1���zS���a���5e'��Ǳ�:���o~i���г���:�/آ�|��&O�9*~ΊR�E2v�G4Y>-��Tv3���K,����Ee�m#<���uUd���^�v2|͖dQ�eb�X����2RE�X2��z��,]��x��\��x�|^y��M拡g['��Ԕv�	�I:�wE)�Mfo�FB���0�d?����(P��K'���G�z>���ӹ1)̻9,M�e���tq���bn~i�o[|w�SwFn�����YT�-����<[/�ѣC�Q�����I3S��>�a��(�y�ޕ'����i�Ԗ:��V�
H�b���W5)QF몔�U�ұ��|�]=����>3F���)��X�e���C9F#F�)RZ�a.��KB�5VMM%�^g��"�������$�j�S�u'(8/�t�#�r}���7�ܳ�.��zg5�S�ԝ�ֻ��ܧ��T�����.�Ȟx������0�>��u'���pl{[�o�(¨��T�
J]aejs\�����ܣ{fDݑ��ˢf]r�ݷcT���NI�f�d�u�9�Q����՛�hh��r]�5\��'6�37ԩ_%8�"��O�^|��ղ��&N�+��S���reJG4�th|)�Sв�O2��78G���"�(Hs-�� 