BZh91AY&SY!�Q �_�Py���������`�z�T(�   `�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L����L���=OH  F� `�1 �&	�!��L�����=CSL&F)��L�=54ޤل��`����~G�	K|�G�B�*$R!	��E1H�.��d��,3�������y����t��T�By~ĥJ�o�t�rq��N.	A��É��b]�	�j����Y���L�z�m661]v-����ܦ,��2��JZ����٘�a�6oRF�m�$5MZ\���ƚ.}��n�͕Y&�R�UWk�]�:)�Q��)ƭ�^����^N�]���l�/�]�i�L"��1�5Ȋ	G�N~s�F&tC�h�dt��4��L�nl�d�,"��MJ/��3�X,��A�3��V��f�
Ջ���2Wz��2�/���$��I{b�,×b�i�'MY�S`��w�ŪN��z�\Lb�:2OЎ#p�""�*���1Lwb7��;x*Mr���e�Qg걂뵰aRD$�3b?���q5��FjD��X�K+[š���@���#QC��,�5�R:(,"$g�J_�i�_�L�k���=�]?�/�����<j�M���	v�w�{���D�h�LZ�b��S�U|��]��������{pmo|pkx�t�|I�a��醃ȩ?H�=(�������&�)�"��Jqsw?b���G�&/oT��ԥ0E1u�G$Y>l�D�:�G��K,�2}��Ec�L�,��o8Ub�͋�^���kY�Q�c�r�-�Q���<p`))�b�٬]���255��⏛�1<$�Z�g/ςQ�}&��qM\Ԧ�4�>
1?gi���C�������zɂ<㽋��9�L%9e%���b9>���tsN�	��rO+b�#�񚹲u�ɵ9T,�K�~�B��k�f͙�Q����d�p�$�Nn�>��$���2yԝ�R:�&�Җ82��F
H�a�ܴ0J�*(�uR��q�X�mQ&�(�w�u��~e2Ff�
`����h�2��F��3f�ܕ%�����-��X�3��G��"�r$�=fuI)�pM�m_b�<{{��>&���Y�H�y�%�S��tN+�;Z��j�=E�{�،דI�Pt{GI8I���s�|��&ֳ���`�7#QKĩ�;T������g��Q�Ͻ��Fƶ$Չ��ǚd]r�կ����zm�1R�g���:0<{�2q���v�����rf�2}j����R�T?��%��`uF�k$r�-�l�tsha;��,iH�eFg�N���-$�(�#Si3�w$S�	 ��