BZh91AY&SY���} �_�Py���������`�      �0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`b`�!�22�M#L&#Bh�4zj7�%w�"�C(��?��-$����d��0��T��,�?Q�1UV��3T�����+,4��x�k���<�]$�xW�*jՅ�-�~kS(�����4]M�]���%�(��gK��)��R�~���n�s)��k6j������\�.�OL�R̯�5W����d����H��Y�C�.�D�s��5��ef��(UUw�E�S�O���"�-��n,:t)i;K��Zd�J˒�eg�`i��ֳ�m$UR]W.�Oz���jk�M�2�7�X�|���ro6�8�h���f����k9M4����Z핳U�3�6�N4�]��p���m�6�*���n���u.VQ�-�s��&Z�Yt�T��O-�y=�R��*�UUUU*��*,��ǃ�j��;�|U)�=VYK���X��a�,�Ҷ��2Ě��0�fl���2���*J�V���kUF)��R)M���M�f�h0Pғ�TvUR�7�m���]_m���]9���u>��j��O�ɫ��|Wnښ�����/��ߛ�T��R�7,Ƀ�N�����]���ɫ�����pqO�96x�t�}���}��I��?�=H����'c{�LاDX~e���)���~�;���2|I�S�tR��)���I�d�4�-���}~�Yg���aIVYf�3�<�.U+%o]b��s���l�)G�FK�[���L��w��%0޳6�af376E��2>1��t,�d�9%��Â}RN���JuI���(�\���;���]b�I���OIy0�8�2}Q��N�ħ2��7ݔG7��a���������o[|wCwFospNu%�Ib�O��S���m4>��8�KI���Q&jtwG��>�%'�f�<�x���BX���RGQ�y��i0��JTQ��)���X��R&�(�y�;��{�f�57�S,�C�-6r��14X�J���	w��ZQ��ji,j򾖱��vǵ�1'�T��+�q�]'���_Sx��Ǚ�,실v�y�u��rN��]��nS�x�$|凙�oF�Ʋ'�Pv����F�����h�6=m��7�GR0�)x�;�z��XYZ��,��:e����(�ّ7dw22虗\�7m��38�'��T���qq),����ū7\��Ry�W}�W03�ͣ����C��N�b�T��>iy�;#V�$s��86i'R�����w�?L�R��1��x�y�ZI�QRF�h���H�
�֯�