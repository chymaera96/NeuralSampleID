BZh91AY&SY$� �_�Py���������`� ���   ��b�LFCC �#��b�LFCC �#S��2  �   S�R  �     �& �4d40	�10T�4�bdhL�SG�Q��x��I�	+�%��3���������d��0TJ�T"�E�'�U�%�d��d��,3����
�����.�׋*f�`�ſ��j`�G%�w|�<���k�g��Ւ�RVnjʸ��K���T�/9^�m���ٶƦ�X.�U�M�.Y��E<�>��6����.�,ٽ�А�6irC|lO
h����ۚ謓D�
����wqԧ�F����s�N�������T���vK�>&~ƚ�JjT��e|��o�n��m��s}�2��=�4�́L*M�e�̯gM�8NJ�e�.��:��XiGH`X'�v���������,�
8�6��l��;y.a�������f�����k�6eL6Yn]��j�cLp����wv�m� ��  �1��,�6����:�}�ڧ�R���>�B붰`�e+I���U>��c�^֪�t��B�*�1_��h��hک��/=M��b��6�o	:jU)F��v��	�c:	2C����7�2<p��@m��e�)v�w�~���͢m4T�-�1`v)�U_?���X��у��z���$��ׁ�O7��k�a��R~�h,yѫȧ�9ڿD���:a�,�ڥ9���Qs�H��/�8*~��)LLE�4��O�;PآXs����K,��}��Ec�L�,����U��5]b��Nv/j��Q�$�n��h�Ix`�RS�2f�v0v��\�ڋ;J>���&���Vs1xN�)G9�0nOt��6t)M�i2{�b.~������ps
3tId��ɂ<�����::�	NE�Ibkv1�����:��l|���mc��::S�rr�eRX�s�r�m_��6g�GW�?5���q��%:i���%/�ʤ�R���6��c�(h�`����M��)J�,إ)��ر�r�5���~�9x>O�L���CS0Ye���xHe#la�X�J����]�f���h�Z�+;�֑��u'��0���IO�p�r����~sQ�6�z�x�GQ圗YNg�Ne�N��>�RG���yZ�5�I�Pu=��8�&���)�3x�OKX�F�*�^%N�ؤ��V�%�<����z�-[j�ě1:ؘ�&E�-M�y�&G���1Zʫ9�
K(�`xx4d晙�y\{�.`2�ɛ��کe7��"��Iy�09�FՒ9&,[�Y�룡���v,>���#�a��*t��Yi'r��677�rE8P�$�