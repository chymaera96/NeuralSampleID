BZh91AY&SY�e�� \_�Py���������`?zK�� �]    SMF���ɦ��4i�4 hSA4"*2dd�F� 2�@��b�LFCC �#	5OU��d4�   ��& �4d40	�10T�	������4d�4z��P��zi���0���$E��Ćr?3�ZH����~�00��.P��-_�IxC%H�����1��:O}nU����I"��]�����e�ߒ����+7��|rrD۝���ty�0$���%R�g
�i(��n�cw�L^�����Jq�ܳ�e23�c��ѵu�M���d�lE��"����`�wP����R���B�x�+e��т݆`6-��4h�����͛e+�$R�W|�t��&��6 Q��X�1C�@a���ʹ�;D-��������o���Ô�����!��4L4�fȇL8�~�к�3�yduG8�.zs-
"�����̈́�J����;�Q[�.Pi6z��|kq��q5��b��S�vG,�%��I`�}�"_���9���X��:�F�lZ�j��2a��Ɗ�$0B�[����=�FJl?0F�n��x�j�A¼����z[��p:�be�d3�����(��5��0ӷm��h�a�P�K{sI�
�g��X��srN3F�C6���H���;���<��t��|p'�la�//��1��IӁ%|�kPjG�1�o��i�w�9���lHB`������;P��c�m�5݊>�lS�R���?U�FK����!Q���L��jIii5d*�f0�2T�Ȕ���(�5��E�Z����Ir�kMhbv�e�C�ġ�'3�D�QT��l�׭{�"��S%���ʨL>��A�QDEXL��QL�:�����=�<�&�EJbԳb��U��Z�E���<�OKՃkrH�F��SȞ_q>��<�H�x�?H�<����'Cc�L�)�"��$S����\�=Q#ԛ�>�*R�"��:i#�,�6��"*:G��K,�2~�Ec�L�,�G�q��l]b��Ά/��d�Q�(E�C��S��b�"��2���fl�.�f����gqG��1>�#a��Y���qޔtS���9�W)�&�'�F"���`�^�{�-�qB�����O1y0G�x1z��N<�	N�Ibl�������S��j{���m��v���tĎ�¤�eRX�s�p�k_��6g�G.��-&NF��2S��${|�IGK���Rw)H�d��T���4j0RG1�<�i$`��JTQ��)��ұ�j��Qt���/��)�30hl0S�X������C)�͚�rT���C4�.�Eb��$b����4��\(���uI)�7��&��.��{����5jΈ�G#�8.�����9�rv5)�:U$}����،׉H��U'�r��"F�����3u6�����̌E/�d�RR�+C��N���8���lkbMX�lLx�E�-MZ�D����6�R������%�r`v�h��33T�<�˽�0D���d�*Cw�NgB�T�?������5���$bŵ���9�G��ذ��Ɣ�	�Tf|i�S�e��%$jm&o�.�p�!��5�