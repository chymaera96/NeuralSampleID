BZh91AY&SYR;� �_�Py���������`_ ��   0`��`ѐ��&��U=OSM����A��4�C@b��& �4d40	�10��T@        0`��`ѐ��&��RB	�dd��M��M2LA���Q������ԛ���$Y$��?��V&��k'�(¢UR�QeI�/U_�It�5H�����2��JO/EqU���ϡt�W��M��Yb���0�<.��m��墱�̔�E%b��z����T�_��:Κ��fv��ͳ�u�G����5i���Zh�r�gڣG-�SW�T3�H6k~$:�ry�U����pr��5R�UW��]�;�����)�]=�
�����2T��:�{��ۤ���KYo�kM������p�.�)�7�rʲ�mR]�e6XJ�Vvae�何WT�M-{e���'f�E>�N-�nZѦyk�)��*ժ��Vs�c�̛��^�`��ژ�-)��!�   &	��=��j��;�}�OY��.���c�ن0��++��of���IU+;Z�}L_�RkR��}�:��"�ڌO���-E�:��;T��6�r��a�%59���|��]H��a� aݿ������,rK�4�S�^o��ScUJdܳ&:���ۋ������s߇��M�g�>�̟K���z�"�X�#{�S�N���=�N�����:�/آ�|���}	�S�tR��)����9���nk"�����R�>L߹�$QYe�H�7��ʫ%o]b���c'����w,d�b��d��<�`RS�4h�va�1ssdY�Q�}S#��Zg['���(�>�	�I:�wE)�&�7�!s�x}������(Q���OYy0�P�d�#��N�ħ2��7ݔG7��0�ꎉ�bn~ni�7��;�9��7k��s�ʤ�m'�s�l�[F�z��4|�7qʑ3S���{|����f�)<T�v�M�bX���RGQ�y'R���J�7]T�9\{�2pP�����^��S4ha��Ye���Z<��3��b4h��%���kD�.�Ud�ђƯC�k]��s������IOK�q��}�����o���~K;"�Ǫs]e:ܓ�:�w<�����>����oF���>������F?����h�86=���7�GR0�)x�<'���XYZ��,�;��:e��onQ��"n��de�3.�jn۱�3��qNՕU�:�\JK(�`��j��44Q�q]�5\��'6�C7ީ?E:���G�O�^}f�ղ��2pl��]�����&T�sLgF�Ɲ�<�ZI�QRF�h��w$S�	e#��