BZh91AY&SY���� �߀Py���������`� ��   �& �4d40	�10���jz�d�ɐbhd i�� �s F	�0M`�L5?UC@ @     �& �4d40	�10T��ђbhji����M=����J�I!�$��L	K|VO��
�UJ�(�������Ipf��f�+,4����WB���<z%��^o56f����E��rY�w���u=gUQu,QIQ�KT��Jp���Y�[���]v9�۝k��9�2�{�vη��sf����l�oT�<3��6k}�$9�d񦫟O���nܬ�R�*����C�O���E6���m/��ٞ1k�&q�3e{2f�LS<�s���e��Sm�EQ��������6�wibn汢��x�d�^��c���,��f�������T-QU&]-�RkQT3R�S���QXWk<tT-�nce]n����v�[֦��iOx�ԙiN@�! �  0K-=g{�j�F;T|�nS�zl��Qg�c���YE����RUJ�֪��ުI�yU�jj���4�bS*�ʑJn��ܻFKA�CjNw�'b�(�@��Ҏ�S�*6�!��L��P�Ҡ(�n��.������[�����7�S&�2`�S���O��lX��Շ���=�s:#���Ο?�O����5E�Z�o|�{���&lS�,?B�ἧK���\�>�'ȝ
�����L��t��O�H���S8��4��ѣ�aIVYf�3��t*�Qf��/�u2y��d�ģ%�;v��Ix��RS�3h�va޳1sf�Y�Q�yfG��ZgK'���(�>sd���)�%)�&�7أ!s�wz�T?���(Rh�%��^L#�<>��S�bbS�vrX���#���0��I�bl��S�޶��<fܙ��.d�IeRX���q�n_��F��Gg�?��f�8Q&jrv�g��I(�yL�u'z���i���c
H�1�Y0��JTQ��JS�ǹc'2�7�E��S�����h��Sy�0��'�Z<L�3��14X�J���	w��ZQ��jhd�����Wg�{^�uI)�pN�'2��I�>�C�oq���uE�;<��t�'bt��w6S�u�H�;z4\�D��T�p�80'�pO����n=m��7�G:0�)x�;�r��XYZ�W,�;b�9e��7�Q���6��de�3.�jm�������	�͒�K:]���;<}Y�f��O;�w��s8�Z<��B�:>Js��"��O�^|��չd�&L����trjbv���R��1��u��Yi'�EI9�����"�(H_��V�