BZh91AY&SY{�Ao �߀Py���������`�      �0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`bc�0L@0	�h�h`b`�!�a4�M#L4)�=F�I�����"[�$X�d5����d���,���
�UJ�(���ת��Ipf��f�+,4��v�W[�xytK���2��XYbߧ�0�;���Z8)�V��W��S�zŲ�
]N��9���Y����gf�:�6h��z�E�\���U=2��&n-/�`Ռ��G�C�6��7��l"��MW=����J�5)B����.�|�na�^덹���g���dњ�=���L���[�nD�2RoR��o�mo6��f�e��ܥ+�O3zח�w,:eXRۗse{��V�Vկ�[���w+]L��;[���L��U���O�^-8^��f�R�Ļ����+���c�ݵ̫��g�3oY2R����Ok�T�)J�ꪪ����J,��ѫ�,�Q�Se=%)K(��Y=k�نYE���-דC+R�2[�TՔ�F�J�֫Z�j�%�eH�6����v�KA�CJN�Nʪ��}&�/w������-t鷷���6�����<��/�v�����.�ix����-�ƪ�ɹfL�s����k�:�5a�v��~N1��M�7�=�>v�=	�����X�#{�Sڝm��0{�����K?�yNnǃ�(��$}�O�8��)L"�<T��O�rƱl���R�?Vo{
H���6��g���U��7��x��d�[,�5fX�q]�d����d))����X�0�Y����,�(�>���7�.���<�g$���u'�$曻�	5����ü���a��\�
M�Y=%��<�������N���bo�(��o�ñ�;����]�o[|wCwc7���N��U%�i?�AO��hѡ������i3v���5;���>�%'�f�<�x���BX���RG�'�	]�EnR��q��d�R&�(�y�:���|Jf�57�S,�Ru���C9F#F�	RZ�a.�4KB�5VMM�5y_cX���;Os�bO�%>�$�$�_z�>g���[��n<Ͻg\]#��΋��7$�Nk�]��zO��Ya�y�Ѣ�'�Pv���r0`���>F����o���1�QKĩ�;Ԕ�����g��Qٗw���F�̉�#���bf]r�ݷ[S3��qN�jS*���Ĥ���'��憊O;�ｪ�q:4yY��Hq���֩��>�y�:�V�$t2d�l�8.�Ʀ's�a�dʔ��������S̲�O*��7:����ܑN$�P[�