BZh91AY&SY���= �߀Py���������`�      �& �4d40	�11�& �4d40	�11�& �4d40	�11�& �4d40	�11�& �4d40	�10T��	��bh�� �Dz�ɦѦ�����Wd�#)!�?�����k'�Q�D��"/%T���U�I/ �R#�H�I&VXiI���\o����붤�3��T��0�ſO���
9,���躛|�,MUj�)r�J����Ժ�R�>r�Vr깜�ߺ��{s��7�dp��5a�6vk;�j��Ʈ����vDp�V$���}���M=����Ԭ�I)B����Wx��>j5�E9���k�����YvY[K�]���FY���]Gf��Ե��D��b�|Z-+�i�����,�k,��ܝ��hT�F�6�*�f��U'<�1ud�z޲Z׻v����гS��uU*C*G�2���k�������&�3b��9���63��c�V�)���a=.�R��*��UUUUUT�%���;_�k�,�Q�TmS�y���Qg걅�ma�,�����F70�{��C/J�kE��RUJŭZZ�_��]�-U"��FS�ڻ6KA�CZNgڜ�U�u&ݫ��o���?ᮜv�z�ta����s�~>Ϣ�i����Ηoix�����z5M���ɱfL�tUW���<�Xz�O[Ն���;k���O���$5I�Š��F�֧�:[��`�E9"��Y��IN�'k�(��$}�d�����)�S!gz�8���lX�"���{�Բϓ7��$QYe�H�9;�z��Y�u���:Y>�ՙJ;�2]bΥ�u�2RE�3��r�,]��v��\�ڋ;J>o��I��t,�d��Ҏ��a�=�N���JsI���Q����<�l?����(T4r���/&�̞����RbS�vrX���#���0��I�bl|S�ܶ��<�L��8����Ib�O��S��~���]����7Q�RI���r{�ǮIGy�3xԝ�R;��kȖ9��V�
H�1��ZJ�*(�uR����dި�t�];�:K��|Jf�57S,�H�kG}��r6�#F��RZ�a.�4KB�5VMM$�cW��5���#�OS�bO�%>�:pCz��I�=�kp��gL]#���+��C�:��wS��O)�T��,;�6�h��Ȟ(����Rs����t��;���9��FE/�d�RR�+S���\]G,������YfG[#.I�u�Sfޖ�fps���Jd�t88�Q����՛�hh�x�{ڮ`g�G���T���ΕH�)��Ϭ������L�7���2�����v,>y2�#�c:4>4��Yi'�EIɣ���"�(Hs�f�