BZh91AY&SY��� "_�Py���������`(�=��   �0L@0	�h�h`ba"��Q�4��4a  2�9�#� �&���0F&���  �     `�1 �&	�!��L���� LL��$� &)�����=Dޤ׀+����3���d	Kw���F
�UJ�%Ģʓ�^��Y%ș*Dzi*I�a�'w_emU����.������X,�o��0`��Λ��L�v���0C��FP0b}{�/TC�׽�ka�̔�N���8�
�Y�W2��,s�]�ر��u�4�sSSW���&�Dӈt�,��$���tA�IBkiӖ�4iN�ҹ��ݜ�mJ�4	JU]O�wi�N�X*�4ײ���˗�kT��]f~����2t,]��y���#.Jf��q��;jRH��	��s�9� r㉍�����r3�*�Ĩ.�e�§��.����I�剃��z\u$]/&�Ԍ����$fH%a���Qу�x��^�����ûvMK$5{�o£ڬ�їF7�Ҿ�R�4�˻�D=�"��
�El���il�d.w��9���p��1R��;$�O%������S�&.+b9��ر�l[��CL��-)��!4   &	&4�e�N������*<ԧ��)e~�D��$�QD!8�Y ���I��S-�%f�����l�ՙ&p̌!�gi�F�H�5Q���.͊�bP�B�|�{M	�a�.8&O��D���=�|~�������b�{�O��v�T���,nK�3�S��<��&�B�1iY��M�U����%�}��'��������*y�D��!�D�;T'��ǡ�E=i�������g��%7���EΙ#�&/mT��T�0E1x�#�,���J���eE,�����RE�93�����U��5��xI���5,�
0eb�i]%I:T�Iu����k2f�v0v,�\�ԋ;
;�9��&��f�7�u�w%���=�M駊��D��Q���:�������(R&n2Y<���Q����8�L%8e%���b8=}.h❆K���6���I�i����bp�K*�ų����cR�ٳf{Tr����9�&Jqt����%'���Rv)H�2MO2X��L��a��Y�
R��4�Jn���bؤ��J.��r�}_R�#3�Y��,��H��h�e!��Q�f�c�*KS	w��ZQ�X���Ƈk��\�B{�	?������l�b��I�|^���4�ϊ�x�G#�8.��ۓ�o]��ҧ��*H���+Z3\M'�*����Bn0�~���3t65����̌E/�T�RR�+A�r·L]Gz~mm*5�1&�N�&<S"떦�\�dmnM����Yj�{kiIe�{Z7��ԉ�m]�h\�e�7k'�R|�s�E"	䗞C�45,��LX�53D�]Z'K�aߋR8&Q�����r�I;TT��������)���D0