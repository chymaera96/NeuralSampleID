BZh91AY&SY�3�� �߀Py���������`� �    s F	�0M`�L54)�z� @     ��b�LFCC �#S�UF�       s F	�0M`�L$ �hd	�z4�Ѡ=FOF�&�n�J�	dFI$~'�`J[��TJ�T"�E�'��S��.�5H�U#5D�Ya�'���+�ww�.����6l,�o��0��w|?T�����J\����y������t�J�Y�e��f�,o,��u�6Ҭdo��o��	�S���ҫK�/���|�S�����m3݂C�5Ol\�?�j�MR�*�����ا�F�"SZ����ZN���ƌ*k뙳���k�2[�ْ�P]I���|���z��T�Sf��c5�ӫ/��ka��-���I�[��٫��*o�њ�WFj��1v�Z�߷gҳa�y�{SeO)�b� ���[AfᨂX(--��-����Zm�ha��t&�ť=� �  �%����~m��e;Uc��OAJii�aK~�I�]v�i��/3���[L��屋�[,�z���Z���am�T�b�F�H�6���5]���`��'��"P ��:H3
P�O�J����㝨��`�ΆO����}�5�6�Wic�.���O��x�Z5M���ɱfL�tUW��k�:yڰ����{㝵��'��'��j<jO�-�J7<�})�������g�ܔ�rw�b���G֙>d��9)Ja�Y�IQd�4z�R*:Y��饖|Y���Ee�m#<��Þ��E��X�?��d�VN�,S8�e����d���Pf))�噴X�0�Y����w�|�I��MŤ�*Y���9s�'��z{d�	����Y�ܣ!s�wz��{��@�CG),���aa����9v&%8�g%���8���Nh��&���F�Gi�6rf�N-�ƅ�Ib�O��S��~����q�֓7a�I&jrv���{$�u<�o2��JGS4��vpհ9�C�9�J�UQE��W=Ǳc)�R&�(�xht�����jn0�Yb�����r���,w�Ija����-��Y54L�5x�[X���;�z�I��$���No_r�>g������x=�:b���q]e:�؝�͊z�I����nF���'�*��{bs�Ls�9��h�om=m��7G20�)x�;�r��XYZ�W,�v��r˷��أsk"l��de�3.�jl���389ӂo��+*����RYGc��Vn������w���q8�xپ�Hp����T��ye�������2d���s.�MLN�r��*R8�3�C�N��-$�#cy4�w$S�	
=0