BZh91AY&SY�y �߀Py���������`      0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��RB&F�'���h�=F�i�m&�"�II2A���~�R���(¢UR�QeI��U_���&j��Fj���)<;{����<�O%e�4x�Ybߧ�ja��v]�~<�y����L)r�J�p�Ժ���Jt}w��깜��uX�7�0��cz�G7�ыlh��f���&��<uj�胚�$�6g�C�6'rl\��;��*�M�UU��Wxε>*5a�^���9o����	�j�S/Lči(�4��l�:�l$�I�YV��b-QJ��Ŕ7�-��)�e���f;�2]n1�F��ś�E5XΓ<9�+��ݕil��lg�;4�Z꒚3��ß�V�*�1ͬά���E9z���Ssf׏�z��)JUmUUUUUURR�OK��5y���>JmS�R���?U�B붰�(��fڒ�V��U�j�'�b��54��U]�E^��ک��1=M���Z�i9�bu)J7Rmڽ��������5Ӗ�W;���i�9�?�����]�m5rv8���^)���O��Si��2lY�j��U���텎�-X{o;ۆ�	�-���<�q>Vd<ƣƧ���ЍϝORt7?4��t���Y��)��w�r���G���'O�ҥ)�S!g��9"��i�xt3��襖|=�)"��,�Fy�5Y(�r�����3j�ԣ�;�,�wt
Ja�fm.��;�f.lmE���d|��A���d�:x���z}RNt�ҥ9��f�(�\�ݦ������(Q��K'���G�x2}Q�'OZbS�vrX���#���a�掔�16>�$�7-�;�gK7�ɽ9QeRX���r�m_��F��G_T{֓7YƑ3S���}�IG��3yT��R<L�k̖8������b	̱��JR��6)Jq��,dޡ7IE��S����)�40��aL,��G�Z:��g#lb4h�ޕ%���KD�.�Ud�ђƯ�k]|�[�����*IO��8D޾��|����7��x=�:"�g�r]e9�S�9�u�[�%I����nF���<�U[�:�L0}���GS{i�n���1�¨��T흪J]aejr\���Qӗg���F��Dّ��˥3.�jl��ՙ��8&�l����w��:�;�5f�(�.�5\��'&�7ҩ%9�
�G�<����j��2omhs.���'c�a�ɕ)�ѡ�S�S�e��5$lo&��.�p� �(�