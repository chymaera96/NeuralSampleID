BZh91AY&SY��Mg �߀Py���������`_z�R�   � �`�2��JMMH�4       9�#� �&���0F&jES�!���h!�	��bhdh�FC�0L@0	�h�h`b`�!24M�ɉ�����'��M6�n$���-FRD�G�~�@���YD��\aZH!C'䲿�%�&j��FjIYa�'�N��~6�%�v��9r�
���.!�(ӱ���zDЬ$�ZF�%�W��n]�կQ�c������Ju�J�,��s9��m����dnX�˅�5LfÁy�]e�i}1��-�Z��/ع�Ǎ�ٽI��Ąѝl�!�0�D�s��{x�o��5I�UU��yN�|Tka�e�n
Y6�:1�>�SEc*��s�kFZ������jƻ6A0��K+�J���Sm��,�tF�&V�����_+�K��4k7��|_��W�$�b�	�D�=KM*X�NsU��a�p��
��weTvkH��Q(��-�(�BB�+�sU�)BWL�0Q(@CN�\b{�%�ul��TRL]iM�2�Q�j�*4�*e4Ui��s:g�j�m{�2�yS�ś���P�;�^��D+@�f��""�EUUT�����Hj�F'�
4�;JlS�)JYE��О��la�Q`���+�,{�KY-e�T3x�23��*�)�Xb2��i�bX���dP�I��$��*�J6�lؽ�\18�-O������$<��LQ���%�N���sK�>�����ԛJ�ɭfL�uUW����e��-L=n�cՆ�>����y����a���	�yU$~Qh,zQ����[k�Lȧ4X~e��l�N�7��(��$}RFO�8*~�jR�E2vRG$Y>*i�i:���饖~m[
H���6��rG��ƫ%m]b��s���lY;Ta��b�EN�d�K<�d))�ՙ�X�0�Y����x|^i��6��EY���9�J:�A���I:�_5)�MS7�FB���0�=��_ۃ�P�M�}��<�œ��9�LJr.�Km�Dr}=���x��s�y�V�ǐ�͛�H�ܜ�ʤ�m'��)�ؿSF�j����-&n��FjswI�I�Q����O)��cЖ8����
H�b)�hL%rR�Y�JS�ǵc&�D��Qt��u�����j6�S,�H��h�g!����ѢǂT��K�mк�Jɨ�H�cS����+�!�H�=f$���S�qN7/�t�#�p{�G�k<^��qt���r]e:�S�u.��kS�;$z���/$j�<�UG�t�8��0}���Gksa�m�a�b7�
���S�w�)u����gk�.��]�{kZ�����#���4̺婯g[T����8&�l����pp),����S7T��P�w�����rh�}J���S{�R*�O�^|���زG)#&M͍!7��mF's�a�ɕ)�ѡ�aO��yTT���J���H�
ɬ�