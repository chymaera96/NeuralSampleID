BZh91AY&SY�3� �߀Py���������`�T@�օ   ��b�LFCC �#D���z!�h��z� h��0`��`ѐ��&��SBiF�P�'�444h M� s F	�0M`�L$@�ddh"zhO��4(����&� ��	i	�#9��-!�������`��T�E�E�'��&��/�R#�H�@���;�:h�����B�QE8���D� �߃��s�#�M�a�EI�lܲk��JW?����p����U�B˹W]��c��A�d�3i2J��'�P�	�k�$��9a��#6�����5.~�������3�(UUu�˼�<f�%7U�����Þ�A��X�+�V1��fӍҞ����f������ceX��2��n�}�vF���6DL4��g���	���l`E�p�֙"��:�r
w�����$|�¥�8�U��^�,��Ъ����6Al䵱��2Q"#(��]�p�x�B�%�I$$�Hd��}�i�bwX���J��kS�zl�K2)X�c�aDh$�؁3�ߌJ���L�p ��0�ӎġ'��&a)��c�vlV�����mR8)J!)�c���u��ͤ�,��1���l�F� �|Wj�M�E��w#;�>/��D�h�E�G,Hp��In�x1��	<�T�9d�f��75�]�������F�Ȩ}b�X��ç�9�T���8"���~͐�3���(��${�ěU>�
R�"��:)#z,�ƥ/U)���C�n(�$C0�Z�]��ў�
�6.�x)���5��J:\V2`�n��	gd
J`س6k`�j̅�Mh����嘞0�ZI����]��G9�0r'�I̚�)NY4�>J1>������ms
#7	,���`�������8qL%7�e%���b7��&X���S�ޞVŶGQ�j����D�R,�K�~�❭k�3f��(���i2q7T�����{��t<�N�'j���I��K�CF�$r�C�9V��V�*��5]T�7\{�1r*I6IEӻC��GЦH�����LYb�����RH�Fl�;R��0`�z٥�u+�p�cG��i\w�0��fEI)�7&�9غO���6���|�s��8��z�)�ܜS�w[R���RG���w�#5ᤉ动8�Ì7C�~���3t��[dp��F
���S�u�)u����rΗT]Gz�6ƥؓV'S	�u�SV�v���ܛS��UYg3kiIeX�Y�sL��#��wɢ�(�ټ���Hm�S�Ω#�O4���Z��#[9���C	��XxbƔ��Tf})�S�e��E$jr7�rE8P��3�