BZh91AY&SY*�}m b߀Py���������`Q ��   0`��`ѐ��&��SD�*x�� F�   0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��RD&FSd�'��24����h�f�m&�+�IdRFr?��XL��O��D��A.��*O�~�*��]��G�����a�'_*ܫ~Ovat��i�F,[��-L(�����f�Εb酹�r��2�6v�!ZQ���ԧW��Ś���dj�civ�k��o���*vZ���&��]��(��Ue1���ĝ�h$lc��	��x�Eϻ��k��3IJU]���㒞
4`���#��ºj�i9K��v
���=ET�1�p^��
_��i�H%�fa ���@@��bM���M��m����rR�4X{�1�2
F�Q��V����D�N�"B��i��b*))kQ;�BMA��h����
0LB�〱`�8�.;a�D`�:�D\�;�zSi)#4F����b�^�b�"~9�U�F���,A#2BMGjX,�G/�vŵ��s��tD�!Kd���UURRK-=I;_�k�sQ�TMjy�E�R�,��`��l`��J�?&(.�Ȱ"� ���3+pqV�fI��wt�����B2�8�d��V��t��ܩ¡TR��kּ�o���/n�o��(e��O&��Ó�A���e��v�w�}����D�h�LZ�b��S���_]��ս����zpmn�|#{[��O7��K�`�w)'��ǡZ�bu6?4���8���Y�6$�K���\�$}�1}	�S�qR���Y⤎�x3�-���}��Ygɓ�`��+rgd�����b�͋�^�u1}Mk1�GZ�WX���'6+Ix��RSř3X��;Vd.jkE��$��$�f�t�x�;Ҏ��`ڞ�'Jj�:$�d�(�\���K���nt���d�yG{�?T��0��]��&˱���:�]�;L&���<��l�g��œē�jp���,[9��
v���͛3أ�\�����I�����=�J<O!�ʤ�R��d��d���4j0RGA�;ӡ`�+����U�JS}Ǳc��%N���|_�#3��0Ye���Z:�He#\a�X�J����]�f���h�Z��cGs�i\�I=oQ���RJ}M�j�I�>�絰{�G{ܳ�.������KzrN�ܝ�Jy���Ia��#5�i"y"�O`�y�L���������z�#�lGB0U�J���IK�,��u���qǟ���Fƶ$Չ͉�Ⱥ婫_SD���rmd�Ubt�7�QɁ��ѓ�ff��.�4\�e�7s'ک�E:J�A�'�/>��4kY#�LX�����š���XxbƔ�	�Tf|i�)޲�N�$jm&o�.�p� U@��