BZh91AY&SYO8% _�Py���������`� �    ��b�LFCC �#T�ڧ覙 h�  ѐ  0`��`ѐ��&��0`��`ѐ��&��0`��`ѐ��&��RBLF�	�i�&���h�b�m&�v�,!H�g�d0%-�Y?�*%U*D\QeI��U_�Ir�Dy��I2��JO��\o�~�h�wW��L�X���Z�aGJ�۾_��
g���U<�0��))��+��n�����)��Wr�s���Ӫ��{F��s�-��l��7SkW�S��lc)��<���I!�l.Ho���.{?���7+4�R�UWk��u��Q���,�VOUC����Z�FyR���WV2������^�͜���d��,���Ѝ�kW�f9�M�g��3i��}�����*�pZ47�-)T�K)T��'%Դ�V�8�jɥh�fL/c%�2��B���F �u�Z�Y"��٠�X��e�|�}��hf�J�i�u��M̖��)\�Ye���75d�=�aQjn�x)�OK�T�)J�ꪪ����JZzs�j��;}�6�yO2�*]E�E�.�k�F
k6ԕR����kUFJG�b˙R٭�S&Z�hҩ�2�ɵR)M�e=-��d�6Ro�P��6�^�eo�m}s����o����6��s�-_���f�j��,qK��^)�~O��Si��2lY�j��U���텎�-X{oKч3�>1ŵ���O���"5�-�27>�=)�����)ҋ�g��)��w?R���G�2}��S�t�Ja�Yޤ�H�}ZDl^��楖|�=�)"��,�Fy��ƫ%n]b��N�O��fIGS+��[��d�"��
Ja�fm.��;�f.lmE��W�d}���h�9�;�O���s'�IΛ:T��5���2?Wi�����ps��2Y<���<c�����=i�NE��bn�(�OOQ�K|t�q���rOrۣ��:Y�Ó�9R,�K�~�B�ͫ�h����ꏊ�f�8�3S��=�c�$���jN�)�i��KY�V�
H�b$޲0��JTQ�r��q�X�s*$�%O�Ax>O�Lѡ���
ae�*G�Z:��g#lb4h�ܕ%���CD�.�Ud��d�����W_!�=OA�?�����S��2��I�=�kp�޳�.��x�%�S��:ӝw[��O)�T��,<Or4\k"xb���u�&��S�h�s6������U�J���IK�,�NK�u;"�:r���6(��ț2;t�e�-M�z��)�9�l��������������CE#����s8��<߂�8}���T�G�|����j��L�ͭ�tt�1;��L�H�΍�;�<K-$�(�#c��?���)��y�(