BZh91AY&SYB�� �_�Py���������` ��   �0L@0	�h�h`ba��bmOBdф4�C&&@@� �`�2��j~�@  �     9�#� �&���0F&
�A42LM	������G�6�v$WlH��H���h������F�����ʓ�^��Y%�5H�M#5"ee����Nj�W����.����3x�Ybߧ�ja�Vv]���y��}L��(�����)��T�?��՜v��fi���s]�ܱ�W��=9�R����>����S6�J��`��͙��捉�M��o�߱��U�k)B����]�:����咨Y�^�\o��2��)����1�服^�x�lFU!���%.�����K�u��#U/�x^D�dnpnp���ʺ���M�]}�g|��%է	Jo��۫fz���0a�x���g�-[����etک2P�2��ɛ%^q���5^�ݵ̭��3j�&2���Ʀ��Jz!A	   	�M2��~��<`��G�M�y�R�Qg�h���k0����l�IU+e�UkZ�֍Mq�dͣ,��zM��Jm���l]�%�ȡ�������(�I�j�}��ꦒ� �,\ʄ����j������Er��9���/����F���R�6,Ƀ�N�����v��O;V�[��a����;k��'���a���G�S�AcЍ�*�Zt�?4��rE�ĳ�n��rw?b���G�2}	�S�rR��)����8���V�,���R�>-k
H���6��s����E��X�?��d�6��g,v�d��x`�RS�3h�vaܳ1scj,�(��s#�7�EY���9s�'�a�=�N���JsI���Q���;L=/l?@�Q���O9y0�0�d��Ꜻ��K����vQ__�Ó�9'q���8���m��xM������QeRX���q�m_��F��G_�?��f�9�D�NN����%O�̤�R���6������RG1�w�2ф�*R��6)Js�{2oT&�(�w�t�����jn0�Yb���r���,w%Ija����-��Y54�,j�>Ʊ��u�[�bO�%<�t��z��I�>���~ý�Y�H�<ӊ�)��N��]��lS�u*H���3r4^k"x���u�s���t��<��9��FE/�l�RR�+S��d]G,�=�͊76�&̎�F\�2떦ͽ-fg:pM��-iVt88�Q����ћ�hh��8.�5\��'�7ةE9�*�Q�'�^yL1�j�fL��ZG2�����v�>Y2�#�c:4>�)޲�O��67�G�rE8P�B��