BZh91AY&SY���> �߀Py���������`z�P5Z�   ��b�LFCC �#	M	)�4�  � ��b�LFCC �#	5)#   �    0`��`ѐ��&��RDdh"zi10����d�����m&�$�넖�1�Fr?C�Z)o�B��*$	d�
=��Y!*Dy�)!���wvv7*ߛ�ݜ��TX�$q���a�$�7p��屑�oB\.�[�,$��6X�	����c�ʷj�L��66�خ�i�c~�f����*��U�S��57ośCΒm�6"F��9`Hm�)ؚW=��f�l��3�R�UW[�]�9)�KS}X�����*��"(��
��T���t�K,"��ӸmX��g8������?��k�"f��VWZ���]RJlm�����iH-�gQ%����q���>"��b�YÂ�ɵtb�&�@��TLYBڝ8����!�dz���ADiyVBz��*VKs�3"�]�f�h(S^�C�t��+=kF�X}N�±,=�ܑ8TF%A�*G��sJ*���l�`�o:bB�%�I%UT����2L�Ը]���0C�I/�vC�㈁�q�H �$��ev�h��T�T�Kφ���l-Ÿ*��Uh�b%2,U�!�Θș�#(%�� ��ġ��k�Aڢ�k�թ{�����z��vw�5�$�>J]��^��E��Xޗlgx���pxfК�
�ťf,�9�����K��=.O�����>Q����O/ğk�<�h%I?X�<���)�';[�LLS�,>���\���.�Ԣ�T��b�r���JSSgE$pE���F����=�jYgћ��IV8��2�I��o��E��X�?���5,Ĕt��u�-]EC�LU$]�B��5�ɚ��,�ڳ!sKR,�(�x�'�I����f.Î����6'�I̚x�M�h�=�1>������ns
n2Y>��`�������y&�����v1�I��lqN�	��pOZ���4�d�plN�Ib����S��~flٞ��c�ZL���$2S��I���%��Iڥ#��jyR��P��`����M�A�S�IF������R�-��k���v���7̦H����`�,�H�����R5F�5�ԩ-L%ކih]F�b�g$�cC���DW.����I��$��ޛ�6/�t�c��������{�s��9��)�ޜ��w'[J�yЩ#�Xw;�њ�M'�*���RM�L��7�������5��0���TR�*uε%.���,�uE�qǫ��ң[Si��bc�2.�ji���$��ޛ�c&*YVs77�QɁٹ���ff�;ۗ{�0D���d��Cw�M�uH�?��K�!���H�$ŋcS86��-�ְ�ō)���Ӡ�r�I<J*H��L��]��BC���