BZh91AY&SY���� �߀Py���������`�       � �`�2��� �`�2��� �`�2��� �`�2��� �`�2��*H@D��14�4�����z�'�=55=�8`+�	`��G�?e�����d��TJ�T���ʓ�^��Ԓ�3T���3T�ee������U�<<sE�Ƽئo3,[��V�Q�g}��G�N:C<W*�LRWCJզ)u<<*����Y��3�����p]�븜2*��/�8�e[��h�1�/�س<��\���$���.$:#d�˟w����ƫ4�R�UW��]�;��(ٶJ�gU{�1(�w�[;��3d����T�:�]��cܿ��K�#�	�����V�:6hϢ���g��Uy_J_nN'�+NM��m�k2�gRe�/k�6l���k���/QZ-0���V��Lpj�U3�j�0�kijn����n��t�nV6�Y�5l��Vy�p�\�n��ݾ8�,ẘ���Q��m&�{^*�)JUqUUUUUURP���<_��,�Q�Su=%)K(��Y��n�,��|�pdkZ/v�������V����UI��KTn���b{[�Ւ�dPړ��	�IT�)7�{����Z���5Ӟ�ާC��7���d���������zj��,t��Z^)�?�7�F����2l�&:�����:�Z��;���.P��Kw��O��'���֍G�C��AcԎ�Oju�?T��v"��Y��:���Qs�H�FO�9*~��)L"�;i#�,�&�kC��~�Ygś�aIVYf�3�y܎���Y�u����['��d�(�1c��w�d����d))���X�0�Y���tY�Q�}#�8)u2yNΔ����8��$�M��D��ߊ�����a�}���NN�B���K'���G�y�>��I�ܘ��]��'�����;؞&&���>��Gy�6�f��S�"ʤ�m'��)��~��b��${֓7q�@�N�x�}G�$����
O)��w֖:Y�V���bt�YJ�*(�e)N���c'$�$�����/��)�40��aL,��H��G���r7�F�<R��0�]�h���j����5y�kX���;���1'�T��K�9Hq_��>g�����lyߊθ�Gq��YN�Jw'R��e='j��Ya�z��Y芨;�`�&��)�4y[���Ќ*�^%O	थ�V�5�<����̻���pnțdw�2�LˮZ�o��frt�$��T�kY���RYGs��Vn�����r]��\��'6�37ک_5:j�H�i�KϨ���Y#�ɓ�v��]�LN����*R9�3�C�NҞu��y�T���4���)����