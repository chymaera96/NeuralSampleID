BZh91AY&SY��
& ߀Py���������`�      �& �4d40	�11�& �4d40	�11�& �4d40	�11�& �4d40	�11�& �4d40	�10T��hM&&�ji����G��&jj{Ro��D�D����?u�����d��TJ�TH�(���W���$�C5H�����ee���^>��U�G��B]=���s6X�����Q�g��/�E����]KRT�-L)��T�/a^u��������ͳ�u�NGܻs�역����jj�jf�a8�;D#s[��!�7'�5\���Uf���*����Aܧ�F�N���{�*L�:VW�{݉;�t�6����&��)��2{gbɗw��)�d��
��[䭩�?���:3i���*]���x���%��ݺ�[9���	��\ɭ��qb��k댴�L�ꯎ�Lh�^����7*4��8g|���p��o�-yk+7?~�7Z՞�ecuK]�^�W���=�R��*�*������)Z{Q���^��gz���l���YeQg���a�,�Ҷ��U�k�m1RUJ��Z���U-��UP�6&j�L��/*E)���˳d�6����vUP��6�{���m}s�Z��ow[��6�����&����]�jj��,rK�4�S��7�F����2nY���uU�|mv��g&�>�s��a��#��<�R}��>��a5�#��Ac؍�Orv7�T��tE��Y��N�G��(��$}���'R���)�S!gm$sE���bZ�I��?e,��f�0��+,�i�'Qʫ%o]b��I���l�(Q�w,fŋ;�)"�<��z�,]��x��\��x�|�T��#yh4U�l�s�$���8'�$�M��5��%�����~��z�b�GI,���a����G�N�ɉNe��bo�(�ow�ã�tOs�sO��m��y���Q��9�,�K�.b�-��hѡ�(��G�i3w�jtw���t����f�)<T�v�M�bX���RG�N+	\ԥE��R��>匜�Qt���/��)�40��aL,��D�����C9F#F�)RZ�a.��KB�5VMM�ƯC�k]��r=�i�?�RJz\��#���I�?S�o���~K;"�Ǫs]e:ܓ�:�w<�����>����oF��Yꊨ;�p�G#��_��>f�3�c��x�qFE/���RR�+S��g|]GL��-��7�dM�쌺&e�-M�v5FgS�u'j�V�u��E%�w0y���u�OS�w��s8��=�z�:��qv*E�'�/>�dj�d�hɓ�f��:51;��&T�sLgF�ʝ�<�ZI�QRF�h��w$S�	
L�`