BZh91AY&SY.��� _�Py���������`��B�   G0`��`ѐ��&��SRbbL�      �& �4d40	�11�& �4d40	�11�& �4d40	�10T����&�����SF�5='��I��-	2�H�g�h�	K|�O��
�UJI�E�'��S��/$3T��R3R��ғ���E~n���]/W�l�Yb���0u�w|?=E,ԵLHiP�����zBv�_Uh��	��JWG���v����[��r��Cr�G.w,��y�2��1�V����_eL��a�Љ��5�v	X�<	����5���Y��)B����]�;��و��U�/')��4�Jd�\�3Gn���cv�z�^��Rh��|rR�����^u��EV��HlUH.pZ:�9�KdK
I�Q�f˩ˮ�e��/}����ܵ��{�cU�1�'�r��(D QϭA3�7*�WK2�_V��[kel�#=V\�ڶ�mZ/��n�"�J���Q(��u��=�lf!!B�$�I$2f9���G�Y����v���M�}e)��F���dz]��d����|�g�bSm1sJ�VX����|1j�^��Ui)jU�LF�H�7Q�17.ђ�`��'�#��	��jP��y]���U�;�(���L�����.�u5t�K�w#K�>������7�S&�2`�S���>�]�c���c��z��p'�9��o*y�},>�y�j<*��E���F��O�:ߢ`�E8���Y�7ȧ;���\�=�2}	�S�qR��)����:Qd��*^�P��gw��Y�f�XRE�Y����p梲Qf��/�:>�哭F��v�n�FJ�Ja�fm.��;�f.l܋;�>o��H�ZI�����2Q�y�9�$�M��NY5���2?gq������s�G,�Yy0�(�{c�N=��N���7ݔGK��0��)�bl�)�o[|v�n,�R:\��Q,�K�~�N����4hz�vu��ZL݇5H3S��G��z�u<Fo*��JGS4��%�fpձ�$r���9V����*��,�JS��ֱ��P7�E�ǩ�^��S4ha��Ye�I�-l�3��14X�J���	w��ZQ��ji#%�^��Evt����ğ�RJ}Nd��Ⱦ��}���o���{�tE�;,�]e9��؜�͔�ΥI����E�k"x��ǬvH�1#���d��:܍ǥ�8���FE/�t�RR�+S�rηl]G�}��ondM�;YqLˮZ�n�k#3��8'#6T�-g;��Ie�Y�憊��p]�j���N��7�R>�r�"�	䗞CDjܲGL��9�D�]Z�����&T�t�3�C�N��5��xTT���j��w$S�	�.�@