BZh91AY&SYpd�� �߀Py���������`�@
N�   `�1 �&	�!��L����i���M   hb  � �`�2��Jz���M=L��     9�#� �&���0F&
�A24��ɉ�����'���M6�vWpK"2Hi#�?E�R�+'�Q�D��B.�YR~k�W��]j��Fj�2��JO7��*ߋ��At�y��՛,[�|��Q�gm��G1�ҩ���%D� �ڬ�LD���\�ks9��U�捭��nX��V)�vǩ�e�[E��V�fjٻ%��q��hHf�Z�!�Ț�}��~�ݵY��JU]��w��S�F�Mj����sԴ��\̙2h�S?b�ŝu�lK��Yj�l�$URZ�|Y����o��9���g�2��a��yҬ�i���es\��VZ���߮M[U~;\�k�t�%�[vݍ��}thҺ`�-�gS_�f�͹�۷6ܭ�d���4�ɭ���V�7є�S���]m�o����q>�yDDE�*���$I1�Fy�[5��,�Q�Q�O��Ye.���c���YE��e^:/v7,̩-��kF%�TB�I��Ғ�(E �bK�m�& � [H�q� �a�YaJ��9U���p�L2D#	P}qcD����R����E8���^)���'��Si��2lY�r��U��-v��G�=�ǭ��{���qmu�	��������*��AcԍϡO�:��`��:Qa�,�ے��{�(��$}i��N
���JS�BΪH�'�bƱ���R�>L�c
H���6��i��q��E��X�?��d��GZ��X�Y�v���.�A����f�b�,ýfb���Y�Q��L��n4]9�<�O����oO|��6t�Ni5��
2?Wq�������2Y>��a������=��NE��bn�(�O��å�)�bl}�I�n[tv�CgK7RroNT,�K�~�B���h��(���i3vi$�N�j|=G�IGS�f�);Ԥu3M�JX���RG1�x'2�	\��E.�R�n=�7��t�]<5:��|Jf�57S,�P�G[9�m�F�;Ҥ�0�]�h���j���&K����Evr��{I�U$���8A�}ˤ��k���>�a��,苤v��u��qN��]��lS�:�$z���.�Ȟh�������`����<Mm��:Cp�s#
���S�w))u����rηl]GN]��sb�ͬ��#���Jf]r�ٷ��fpqN	����T�pp),������7<��C����s8��<��Z�8|��t*E�>�y�:#VՒ9&L��Ze�����w,<reJG$�th|i�S�e��U$lo&��.�p� ��a2