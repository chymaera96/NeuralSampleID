BZh91AY&SY9��� ߀Py���������`�@�&    s F	�0M`�L%L��)�d 4     ��b�LFCC �#	M!�~���d   h  0`��`ѐ��&��RBL�@�'���MM�=F�I��&�nąwDKBL�F�?����)o��(¢UR�E�QeI�?DŪ���"=T�ԃ+,4��������t�_���ae�ߒ��
:u���tx)��f,��T0@�S����JwQ`��ϼZ�7�U��r�s9��[ˮ޺��s\���w�y©�e�g�+��Uu3�\��]�ԉ��"3k���byb���5�ݵY��)B������x���Jl�����F�:q&��1�f�[�۰�v�7��
�Q��m�U9��/ko�����Aq]�Te�VH-�
��\���X,�!�'%
�)i�JBv��-�"[��TFI��$+�N���n��Z��6)JZ(��-"Td��F*+΢BQ��Ǌ@VD[%2���SE��G"�6�|HB����BI$�LÎ�L��ԩ�����U���T��SK2�)c�h���ma��.��9l4��Z��ؾ��[!�5Z�Ʌ��l�T��(��]xک��>�&��2Z5����j�R�ܐ�H�ėq�f߄�"�wˎ*�}�Ó���f�j��,s���/��ߋ�F���R�6,Ƀ�N���|-v��O;V�c�����O�s���t�{���!艨�G��ǥ�J�Zt�?$��E9"��Y��H�C����\�>�>d���)Ja�Y�IQd�h-�e�J�GK8��4�ϓ7�(��ͤg��z+%n]b��ΖO��d�Q�r,Zv����w��%0ܳ6�af�366����d|�n-$�RΆO!˝(�=��t&�JS|���������������*&�RY>��aq����9v&%8�g%���8���M��;�M�{�y������ɛ�G2q��U%�i?gN���4h{vu�ⴙ�z�f�'l�w��I(�y��u'z���i��K��a�$o1޴L%8��Y�J�s�{2s*�(�xht������jn0�Yb������r6�#F��RZ�a.��KB�5VMM$d����Z�Wg�#�z�I�U$���N	��]'������6rΘ�Ga�WYN�:v'B��sb�Qԩ#�Xx<���yȞh�����9�H��?c�<Mnf����p�oFE/�t�RR�+S��nغ�Yv��nmdM����&e�-M�zZ����N	��L���C��Ie�NY�&����p]�j���N-Vo�R>jot�ED��闟I��5mY#���9�ZD޺951;]��R��1�u�Yi'�EI����ܑN$~!��