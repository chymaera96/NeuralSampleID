BZh91AY&SY��t �_�Py���������`� �    9�#� �&���0F&����$� � h   `�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L����LM4OS	�@�4���4M��Ē����I$��Z	K|O��
�UJD^J,�?꘵U�yj�5#5$�Ya�'���+�w�g���͛,[��֦Q�ge���E���sE/S
\����N�b���+�����\�fl����.�I���F[�R��ާ�p�z�d�)�}�䩻��|�!�Đь������l\���I)B����y��>
5��N5ּ|�G*Xu�ъ�%M&j1��h�����M�%Ԛ(��z�)���7^���s�<8߁���u��\tk�>j��k��y��*��i{�[0�v�S[gn��UZi�Xϥf���!�b��q���)��-�h$�Ţ#j���v6�iO-��\t_��ǂ�JR�\j���UUT�%���<�{�,�r�|U&�OI��m3����豚붰ƙ.��r�O��{+�e�5Z�/����ʪ��Z�x�E��i6�E)��cj�Y-
)?��Ϊ��&�v�w�\>�_\�v�s����}q���L�ϋW���Wl�M\�Ŏ)v���}o���Ѫm5T�M�2`�S�U~~�]���ūc��{p��=�ŵ���'��퇢�*��b�X�#s�S؝-��0|�N�X~e��t���x?b���G�&O�8*~Υ)L"�:�#�,���Z��Tt����K,�پ��Ee�m#<��p�Ed��ˬ^�t�|��2�;X��,�(ùd���d))�r��,]��x,�\�ڋ<
>4��ɸ��EK92y�)GI�0ޟT��l�R�k3}�2?gy�������9
RY=%��<�œ��:�S�˳���vQ����Du'����9���m��y�L�rsoNu*�Ŵ�����j��4h{Tv�Gങ�N5$�������%o1�Τ�R���6�	c�8j�aI!�C	\Ԫ�(�uR��q�X�oQ&�(�x�t������jn0�Yb�����3��14X�J���	w��ZQ��ji&K����Ev��|�Y�?����S��ܺO���>���س�.��y�5�S��v�%ݮ��='Z�����yۑ��k"y��״v��Ę>��qO�������GPn��aTR�*w��%.���9�Y��˻��أsk"l��deԙ�\�6m�k&g���j�ʪrpp),������7)����p]�5\��'6�+7Щ:*�P�嗟)��5mY#��2omi������w�>2�#�c:4=��)��O*��67�G�rE8P���t