BZh91AY&SYn�H� �߀Py���������`_	U��    � �`�2��j`F�T � �4   � �`�2��JhA4�!d����  � `�1 �&	�!��L����LL��OM �=L��S=MM�MW�%u@Z$�$����~�@�J[�d��/TJ�R$�H�ʓ����UZHLU"=4�T�0��*N�}4W���V��F�T�#���H�xs�o��A�T��"���dM;5C����kr��G����eV�ew4 ���M ��q��#q4��*:q�Bz�)��5ce�,v�`у7$&L��y!��4.=��=�U�e$R�UWS�\�8��%�)���g'C���ͪ�VdIQp";�s�P�Ƴ��2��bDf!�&q1��+�c�ԉ�'9s��m2*�H�\EY<���Xh�Zj�$�m@��eq��A�P}�E��byt*T=D4����I�w:����(p�Z#L;��A�؉V�
���_U$W%�d؃(j/k��+�2%�X��AS/}��vJak�Y��
K"�hh�q*_!S�LO7)�HB����R������-=RGc����ye9*ǉ`Gh78�ܫ�'�q��`�mB�g�l�I�>Be6NÉ�M�DB(;��M��h��:dQD	�q����=l&��X-��?�أ� �͚̄l`�<O+���/nr�&$�>;�?��o��⹣M3or,mK��]�����K����2�!�#y%��x2���;�/[�{[`��mit����'���4&c�RG�-�B5<�zӝ��K�dS�,?B��H��c�Qq�H�I<I�S��)z)����7����-M
YRU�c�襖~�^��H���Q�2Gsf�+j\�t?��`��V`�:T`��,�W"���%θ1���f,�.^��b�EƆ�Y�Q��L#Qi&J�n`�8mJ9�1{Z|$��G)�&s�F���/z_��P�L�$�yˤ�㹃��p��o.c%���޾��4pN����oO#Rڣ��h���$okM�	eRX�S�o�i]��&G�G��+I�������������(�y]�N�)SK̖6��m�H�/�rs-	zV�*��4\�R�nՌ�5IE�ݙ�]��)�2/fj/R��X�O�t���F��2d�ؕ%�z���d���3V̤�3v���+���H�=E�~*�S�mM�5�Թ'��l|���w>K9��'|޹e76�ܹ��Ч��T��,;��H�t���䊨8������H��߹�<�-m'��8�|s"�QK�T�JJ\���7�,�r��p×��УSKh���Âb\��4i�g$blmM�����-T���RYG�^�l[�FJ��l\�3\^1�����ܩ�*s9�"�?��˧����VH�$`����'2�pf_9:�0�#z_�Jt�Yi'j��45�'�rE8P�n�H�