BZh91AY&SY���3 �_�Py���������`_U��   �0L@0	�h�h`ba���2�Ph       9�#� �&���0F&� BiMPh44    9�#� �&���0F&
��224L�����jh��'�OQ6�n+��Y$2Bi#�?E�0%-��TJ�TD�YR~K�W�$�H�R#�H�P���ғ���U~��ȺwW~)����-����Q�ge��E�iiA�L6Te!u�U�qB���.�Ȱ�ے����r��Xj0I&��&	q6R�8���fL�e�k]����$s5e��<kO"k\�?�6�h��D)B����.�9)�[�%P�}q_�[ʮ�^��u���,�t��ˊik:�o�`���=��P_H��H�h�H*�����"G��̓Em!�g��u�Kj�c#1֮�lq��޹���DjRVy�'LW�6$_�iU��!n��
W�.R�L��̀�걆W6qC�]"���I3��T	I ��vhqP�41<�I	��j:)T(�1�NW4����u��E�qQ�nl-`o��kQ�6�X���id^\S�LR��pG!��!-�UUUUUT�����;����v(��l���,�u~�A��la�,��8�\�4Q	Bɵ[M(҈���E��`a%-rJ�b��rYA��#4���v���"��Nw�N�%RR���3&NU�����|�槂
�߾T�o>��L���acz]���O��x<tjM��Jdֳ&�:*�����;ژzܞ׫f��olu���������#P�R�Z�m}*}I�������g�څ:]�آ�d��C'̛�?g)L"�:�#�,�-"5��q��ie�&���$QYe�H�4<��Y(�j����,�Cb̨�eb��X�Y]�H�d�E�H3��j��,]��w,�\�؋;�<^Y��Cih4U��C�����s'�IК��Ny5L��������C��΁B���K'���G�x2{��N<������vQWY�<qN�[�pO+j�c����u!�̜(�*�Ŵ����sb�4=�9u��i3r7�#58���Od������Rw)H�f�t���55�RG9�x':�a+����]�JS}Ǳc)̩!�J.����|_��CF�
ae�*#�-l�3��14X�J���	w��ZQ�Y5!�Ƨ{��\�H}oY�?�����tI̾��|ϵ��my��{�t��9i�u��oNIл���OAԩ#�Xx<ͨ�t5H�X����9!��>��oOG[������1�¨��T흪J]aej8.Y�싨�g���F��Dב��ˊf]r�׳�����9�l��Y���RYG&&�n�����7.��.`g�G{7�R�js�U"��闟I��56,���9�κ8���Շ�L�H��΍�:�x,���EI�����ܑN$)f<��