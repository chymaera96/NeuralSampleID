BZh91AY&SY�x� �߀Py���������`_ �]    s F	�0M`�L5CPz��F��4��i� �0`��`ѐ��&��OQ��i�4i�4� �M s F	�0M`�L$@�#FF���4�Ѡ��h�i�m&�"�II1A���~�)o����`��T���YR~K�W�$�I��G����1��:N�5R��v�d];�Å2xX,�o��0`���˾_�k����]KRT�,��N�ʥ7�
�YÅ̦F|ln5`�uۍV1*���nq����3d�hY��b��46Z$�c�C�6'�6.}��v���h�
�����rS�c�P�e]���U���˗�#7[<�d�b�X���ʺ_F^�]M��H`��ܥ��n��7)l�ׁ�L��vs�M[���R�'v��R�$:t*V=�YD��Ti�$�dO&�b�C.V�kf.�^�ltR��D2�F�^�M���!B
�   �����~mx���G�M�y�R�(��X���kQb���Չ�f���H�q`f!����!�[h�z�h�h1(iI��I�JQ�!�@tSq"����J�0��2#���v�(�yAM����Xޗngx���8>��M���űf,�:*����;�0{��ǯ�<����[ʞo��[�cA�S�AcЍ^E=i���&�)�2�᪝.��Qs�H�1}IΩ�8�J`�b,ꤎ�}4���eo��Y�d�)"����Y;����TY�����,^6Փ��ck�ة"�
J`�fl�.�f��QgqG�☟V�k�gC��(�<���t&�*S�M&O��E���`����?�;�P�7,�r�`�(�b���y&������b8=}f.h��c�pOU����l����ܜ(��,[9��
w6��͛3ڣ�\|V�'#}"d�c��=�J:�#'�Iܥ#��my���PѰ�I��Ne��)J�,إ)��ڱ�r��J.��%��>E2FfL�e�*?����C)c͚�rT���S4�.�Eb�͊Ə��"�p�Ǩ�O�%<m��r����}�w���͇{೦.������CzrN�ܝ��yΥI�ý�j��i"x��Oh��`�����>�n�����8���F
���S�v�)u����rηd]G{>-[j�ě1;��L��Z�6��ds��:ndS���s��QɁ��h��33Q�s��4\�e�7��ܩ��ΕH��O$��1�j��nmfs.�-'c�a�ō)���S��z�I<**H��L��]��BB���@