BZh91AY&SY�xv� �߀Py���������`� �    9�#� �&���0F&��O�@       � �`�2��� �`�2��� �`�2��*HA&D��L)�@��D�MؒWl�#)!���|��R�5��(¢UR���*O��&-Uh^A��G�H�I&VXiI���E~n���t�_���ae�~���s������ǜj�,�\���e�ώL�aN��R�<�v���s9���.���p�K���u�S�Ɍ����T�ͱ�ZGn�$4c-�$8F��M�����ƛ�Md�
����w��S�c)�V�Wzë�,8Y/T��3ul;/�i�M�%ԘQe�;h�_�}�p�}�p�+�{�j��67�fb��[%�[=m��e�R�6p�]�שϞ.Ҷl�n�z�4�Yf��SLJ��t�Ai������@#G���P��L
�30��Y��e�^��_5��ӆ}����JR���UUT�����,��I��[^h�e;c�6��<�Y��������c5�ma�2]E�尔�|�/���Vw�j_���a|V�Ux�0�ţj�R�h��6�ђ�`����N*���)Rn��j�{+��k���N[}<�ta���;'��j���E�6�W'ac�.���Os��|�j�MU)�b̘;T窯��k�:9����ޗ��#��f�SȞ_��K�Xj<
��Ac΍����n~����E�ĳ�n���s�(��$}�d�����R��)���I�d��]P�:ǻ�K,��{RE�Y������Ed��ˬ^�t2}M�2�:�k��gaQ��,���IL7,Ѣ��Y�r��͍������̏���I4T����t�%��z{d�鳥Jp�Y�ޣ!s�v�}ol>�ˋ�P�h���/&�&Ol~��֘��]��&번���t�GJw�s�x[���|���ޓ�zr�YT�-���;�W�hѡ�Q����f�9�I3S��'��z�w�7�Iܥ#��6��c��5l0��!�NC	\���(�uR����dި�t�]<Z���>3F���)��X�}�GS9�m�F�;���0�]�h���j���I�Ư�k]|�\���ğ�RJ}Nd���.��{�^���޳�.��y'%�S�̝iλ��ا��*H���܍�Y�Pu�c�Nc`�_�̟3GS{i�n���1�QKĩ�;T������gS�.��.����F��Dّ��˥3.�jl���L�.d�ٲ��kS��Ĥ�������CEC����s8��<�b�8���T���9y�0tF��$r�&M�!�tt�1;��L�H�΍�;�<K-$�(�#cy4�w$S�		'�n 