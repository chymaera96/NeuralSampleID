BZh91AY&SY�|�& ߀Py���������`zPA�T   9�#� �&���0F&	� �     9�#� �&���0F&��D�P4�  �    `�1 �&	�!��L����!���D�0&F��4���lSM��+�@��e	4�����	I|#�B�*!��$1������L�"=4��+,4��������i"]1X��G���-�|V�Q�gm��F��Z��k�X��ɬZH�Ȫbտ��N��:}x�r깜�����z�9�22�r͍�ZeY�g���5�{Z��UbՎ�͎.����VB&��[���&��w��V���4��
����w��S�k����u1)d�u�Y�ߙvj�+-�R�L����i�l�wvvs!3Rj�*��$ݎ{�[-��U&��	_�h	k��
�IK�2�0�TW��ҷZ7����kR��i�ڶ�j⬖s�Psj��Z�U�Bĭj�"�Hw��SC�IZ��
f�C5HU�q� �LA !����\�2Z�B�H���
�А���$
a�ⷥ�0�-���Y�GwQ�92���bct���3s.n�*aηY��L*nSB����g�"".(���U%BYi��~��<`��G�M�y�R�(��'�uۘa��ZU�
����b�eeR,�m-��,�ٔ�IU+9Ie),Qf��h���H�ZL���6Rs����EQJ5�ݹ{����JvW�Yr��/�-N��G&1a��L�jX_3�����{��|�lM��Jdڳ&�:*����K<yݏ;�Ù���o*y�},?y�M�ƨO��ǡ��>��j������g���N��Qs�H�a2}	�S�rR��)����8���V�M�,���R�>,�s
H���6��p��
��Y����,�Sr���Xɠ�,�WiD�BY�!IL5Y�E�������[�gyG��HMMBΆO˂Q�y�9��$�M���<�&or�����a�{a��-�B�M��y�ɄyG�'�?�r�LJq.�K[����:�99�w��_��y��v�#o&n�N.d�R%�Ib�O��S��~����q�ZL݇
�f�'l'��{$�u<�o*��JGS4��%�ᱴ9�C�9֑0��JTQf�)NŌ�ʒF�Qt��t�����l50�Yb�?%����r7F#F��RZ�a.�4KB�6+&�HL�6<o��"�8��O[�bO�%>��C�}WI�>�����M��ܳ�.��yg�S��;�wc��O9ԩ#�Xx<�Q��$O$UA���N!0~���3G[���5�A��s�
���S�w))u����g[�.��]����5ndM����&e�-M��[!37�&��f�d���oo),���Ž���hh��޻�ع��N-6o�R��s�U"�O�>�y��:ccr�a2d�ni"s��M�'k�a�ɕ)Sѡ�QO��x�T���M�w$S�	�ʢ`