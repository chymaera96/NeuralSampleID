BZh91AY&SYI�: �߀Py���������` {@   ��b�LFCC �#T�jz&� Ѧ�12 �2U?F��=M� 4 �@  ��T�  h      s F	�0M`�L$ �&FQ�"i�@M4���m&���"�2!���~�$����d��0��T�!r�*O�z���K�5H�]#5H�Ya�'��¸�ߋ��it��~jd�ſ?�ja��w]��tqS��եWUL��E%u�u��&��S����gs9�����WR�8R�dr�r�6�Jbg}\�8�~&��cF����p��86�lQ�w��ϣ�uqumU�jR�UW����{�na�����ڇl�ʝ��3aSOd��=���5�.��*��3w�u:��84ɞ][������Y����<Y����4���.�Ѧ�k����7k���M{�Q�����i��}�9V�p�"�]�hڂ djSa	)hM���lP��	!��kSRe��!A	   	�M&�e&ߛg�0Yܣੴ���,���Y��]v�.���ѽ�-�vf��f�^ijĵIU++Z�ֵT��6T�Sj1>V�ڲZ��u?�vR�J7�m��}�ꦒ� �,\ʄ����j������Er��9%�^)�>�o~�ScUJdܳ&"�uU�}��qc��V+��{0��|rl�	�}��X}��Q�Q�E���F�Ƨʝ���0{b�a��:�آ�t��>��:)Ja�Y⤎h�{ۖ5���gW��Y�3})"��,�Fy�w�VJ,޺�����O��̨�K����������RS�3h�va�1ssdY�Q�y�G��h�u�w�9%��a�>�'Zn�:��f��d.~�!������8��
M$�zKɄz�����;S�˳���vQ�/�ã�:'��������m��w��3x�n	Βʤ�m'��)��~��2��~I���D����}~��Q�y�ޅ'���4��%�L�q�$u��:�L%sR�n\�9\|�N
��%O>�ax=�qLѡ���
ae�*O�x��g#h�h�c�*KS%�Ɖh]F�ɩ��Ư+�k]��i�{I��$���d�޺O��8������;�Y�H�=��)�䝩ֻ��nS�x�$z�;�ލ5�<�Uk��#�����h�6=���7�GR0�)x�<�Ȥ��V�5�<n躎�w}���7�dM�̌�&e�-M�v538�'�32U��qq),�����Fn�������j���NmVo�R~
u;"��O�^|f�ղ�̙86h�K��S��X{�eJG4�th{��)�Yi'�EI�	����"�(H$� �