BZh91AY&SY�P�� _�Py���������`� �     � �`�2������z��    22   � �`�2��j����        �0L@0	�h�h`b`�!�24L@L&���G��6�~ ��	i	�#I��-!�)o����aQ*�D�*O�z��d��f��f�ee���N���~/�IL�ŝ4xXYbߟ�0K;n��:6So6�j�X�KRV|mќ�8��L)��T�/A]�������k���K�ɾ��dp�r�4�Jz%��E[��XU:�e�6�zD�5�F�].HsƉ�MW>�����Ud�B�*���%��O��E8ײ���,��J���f�3�O�5)�S�k\��ԙ�ʻ�:˺�mI�Q[gt��γ�j���a�P�M�l�\�ɴ䫬���L��αG5�ݍV�vkVR�D4G��RI 1X���rhX,&&�3-2�+J�3/f�>�c���o��h�ͥ��6�L�>bMZS�!BH   R�e�����v��)�O9JQe|�G�u�0�(��V�j�b�����w3g��Z�Q},Z�RfԺ٪�͢��ekFʑJmE筹v�KA�Cu';�'Z�J7�m��}���Z����Ӗ޾�;�mO������~?g�v�����.�ix���r|�j��S&�0w)�U_���n,t�j��v=�f��G��ʞo��K�i�
��E���F�ԧ�:[ߒ`�E:�a��C��~�;d��>���:��0�d,뤎H�|�-RnQ,:Yǿ�K,����Ee�m#<��p8�d���^�t�x�,��)��n���Q���;�f))���4X�0�,�\��x
>o��Cyh4U���Q�y�9��$�M�JS�Mfo�FB���0�����@�R4uId��#'�?T��LJr.�K}�Drz��Nx�O����'��m��w��L�p��NU"ʤ�m'��)�l�CF�j���|�7aƠf�S�o���(�x��U'�JG[4��KY�V�
H�1"s�#	\��EnR�\n=�ʉ7�E�ɡ�^��S4ha��Ye�'�Z;��3��b4h��J���	w��ZQ��ji�5x_[X���;!�z�I��$���8̾��}{���>�q�}�:b���r]e:S�:v;���j�=%���oF��Y�Pv=��LC���)�4w�͏S|u��FE/�t�RR�+S���l]GV]����2&��F]I�u�Sv�-a���8'1�%Jt88�Q����՛�hh�W�kU��rh�}j���S�ҩ#�O�^}F�ղ���'3f�9�GSS�ܰ�dʔ�I����Ӭ��e��$nsG�rE8P��P��