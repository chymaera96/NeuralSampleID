BZh91AY&SY�.� �߀Py���������`�z�U�T�   �0L@0	�h�h`ba�� I��   �    � �`�2��I��jM=5=M�� ��4 � �`�2��*H��i4OBb4i�4z��3SM����ȌR���`�J[�~�.0��X�P��,��Ib��G����Ll�Γǧ}pU����f.��|ir�
����.!���c�牤M<9�g&\H�MY�nff�6lQ5�A�,۝̦F�ln5j�uؚ�bo�r��i)�/�Ec{�v4,�Y�z�7�u�!��;��D�&��_�׃v�d�%(v�����CAr	��,�{�Ro��]�L��5��>ۺe6����K�.4<� d��&��736�Aj��U�7�\j�����u�\��g�������B�u��!�@("R��8x�-*�ֳV��fU����Y��XV2�[-e��\V5����C}6Kpwhφ�m��p
"".પ��%;��9�N�`Y�G�Sj�9��]E��ɂ붮^�TQ�4�,���mT�48�,RhZ�Z�_&k���i6�E)��g�ػ&+A�Ce&��']*�(֓n�� #��e��Z��ۃ� p��"��}iܝR����'�6���R��,ŁާUU~]���ţ���^��$�G�kО���+����?(�=H��S�N���0>��4X~e��T�S����\�$}I��N
������"��H�'Ŝ6(��[(�=T��͓�`��+rgd�.�TY����l_3j�h�Q��-б���y �RS�2f�v0x,�\�ڋ<
>/4��&���Vu1y|R���`ܞ�'Rl�7ɤ��Q�������Ã�P����O���#�<X���S�ra)Ȼ),Mn�#���0so�i�a6>�$�5[X�y��;�rr�eRX�s�r�m_��6g�Gwl~I���I&JstO���(�y���'����I��KYCF�$o0��oX`��JTQ��R��{V1nQ&�Qt���/��Jd���)��,T?����C)c͚ǂT���c4�.�Eb��1X��}M"+���O��0���IO��8A�}WI�>�������޳�.��z'%�S��;��ws��O��T��,<^���t�D�ET�h�N&	����>&n�����9��ތE/�|�RR�+C�坮�u���jأV�$ىщ�4Ⱥ婳o[D���s&+YUgS��Ie�'��S35C��{E�Q93yY>�Hp�)�֩?t���9��6���1b���o]�N����R9&Q��Ӱ���I<�*H��L��]��BC����