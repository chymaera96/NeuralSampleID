BZh91AY&SY�G�� %߀Py���������`yP���    ��b�LFCC �#2#T      �& �4d40	�10�Q)�@��� h�& �4d40	�10T��	��bd�i�i�4h��='�i䛰��H,��"M$��	J�(��"�	%��P��-_̒�	���u!��MTP$�u��_���̒��]��n�X����L0���˾���3����;��0$lS!�C�qm�Y��S���N�1^�7\�fi�c���E�o7,dU�4o��gT�y�f�b�^�����{-m֬^�M�l�My���h�����4mO
l\���m��՚j�JU]����O���9*��5��b��\�u�����d�%rc;�����3�e�����]�Y�R���i���z/H���pi�X��EVS2���!z͔�1HN�T9��Xfe@���:��l%x[�:��V���J����CclũU�[�Ѥ̬�bĲ��T[+4�"k���W��w��E龢h�ҩ��ٶ̷-�9��2L�� =J� BQ��4�t�8K���p�I�
�����A���!4�.r��e�̕"�����ƙ��ضv���U���*���HJ*w�M��m���U6��)JYE�%�<����P)G*hl�&Ad���bS
�]K�]-k]�T�DFA)����M��Jm��ػFKA�CZNg�xjB�n�۵{�u������k����3�m���d�<�_���f�j��,s���^)�n/��Si��2lY�j�U���텎�v�<�����{���vׁ�O/�O�����QޤO�-�27>�=)���S���g�܉N�'s�(��$~�>���9)Ja�Y�IQd��,�"��g�5,����aIVYf�3���s�d��ˬ^��d�VO�3D�c���T�%	w��%0ܳ6�af�366��⏛�2>����:<'.t����7��IЛ9)Ni5���2?gi��쇿���(Q&�RY<���<���������K����vQ^��'4rN�c�qOrۣ��93u"qoN4IeRX����)�ڿCF�R��{֓7Y�HL���D�y�T������Rw)H�f�_rX�g[)#��<i̱&��J�,إ)�q�XɽA7IE�ǩ�^��S4ha��Ye��?���g!����Ѣ�rT��K�к�U�SDL�5w����u�}�A�?5I)�9ӄCz��I�=�cp�����Y�H�<���)��N��]��lS�u*H�7��.���⊨:ޡ։�a����4x�OCtr�̌*�^%N�ڤ��V��<Ⱥ�Yv{ۛnmdM����&e�-M�zZ�fps���T�kY���RYG[��Vn����<���W03�ţ���T���ΕH�O�>�y��:cVՒ8�dɽ��'2�����v�>Y2�#�c:4>�)�Yi'z��67�G�rE8P��G��