BZh91AY&SY�� '߀Py���������`�Ba�   0`��`ѐ��&��P&���� i�   0`��`ѐ��&��T�U@� @     ��b�LFCC �#I@�d��h�SG�h�=z���qv�KHL�H��贆��VO��
�UJ$^YR~K�W�$�C5H�U#5+,4���������"��}4w��ſ?���
8�����إy��Ly��LRVygvuk�52S���N�I^E��ng37m�����]vF匋mpc�A� ��23�]�ܱC��Q'h'42�ѝl�!�O"h���ݼJ�g
P���~��ε<Tja�_]�W,�]:K�v�T���\�׈��{ٕ���
M�-��Y�v��Nj6Ԉ�cb�R��V[��(l��CiQr[c�o$q�ZՍU3q�]���!U��L
�h���_J����AO����ӗl�l�4��hmIx��.�}l����0�;��c��FK��R��ME�����0�Pc��b5&�)��!4   &��-=p�~ng�0Yأ��=)K(��ZOR�0�(����:2^�͵%T��j��{UI1��4^�-Z�͛E��1��b�R�(�}Mk�d�5�s!8�@QCE�w8�g���1}���6�AJ{�M���s4��87��9^��F��jT�Mk2`�S���_]���������=�noG�86:�d������瑨w��Z�m}*}I�������g��
s�;��E��#�O�7�~�JR�E2t�GY<ZDk^�����>Mk
H���6��p�o8Ud�ͫ�^����6,�J0�,Z,v;,�w��%0ڳ6�af�35�"���d|ᴴ*�vO!˂Q�y�7'�IΚ�)Ni5L�����������7��
����OAy0�0�d��Ꜻ��K����vQ_WQ�'4rN�[��Vն�a�5�f���R,�K�~�"�͋�h��(�������59;!����%/)�̤�R���6<�c�8jk0��c�Ne�a+�����j)��ر�r��l�]<4:��|Jf�5L)��X������r6F#F��RZ�a.��KB�5+&�Hd�����+���������IO��7��}����s{��=���Y�H�<ӊ�)���iλ��֧��T��,<f�h�5H�X����p�b>��pOGSsa�m�A�b9��QKĩ�;T�����q\���Q�.σkZ�����#���$̺婯gCT37�&���L���oo),���ɽ���hh�f�����qh�f�!��3�R*G�L��L��d�0ɓscIˣ�Q���Xx�ʔ�)����Ӥ���I;�T����?���)�}��