BZh91AY&SY�$H� A߀Py���������`�zPY+@   `�1 �&	�!��L������ELi4  @   �0L@0	�h�h`ba&��4 4      `�1 �&	�!��L����M�S&&F��=A����==SM��ߑܑ,I3$k#�����P�b"�$�B!A�Ъ�2J��Dz��A��Rw�|��V��/&�.��>Zjͅ�-�>kS(⳶���y�ۊ���j�%��F�%��ái��uR�>��K5��s3�e��m���nX����m�Kl�)��}+Uz��Q�f��f�H���i�֮HsF��&��w�߽ÙY���
�����v)�c�Eu������*�bN�L['1|Mh��eV�V�޹��"��5�5�ITaIk-�fr݆�e��Sb��h�k-��'��M�i�V�$�k/����#�*���R1�
�R�FQ�]�*�XJO���(�Z�IB��=�vKuRA!C��n�2�)'B�"C�"�ZIy�ŬTr�˚��h�M�6�l���_�ݩaKr��S=�x&ќ(�������D%
M��ǩ�kB���!�-�}g��)u~�C���YE�o�7*2^��f[U�kbͭ�ͷ-2,kJ5)Z�e�%��D��fѵv�KA�CZNg�ʊ�J7Rmڻ���Y�C����p�T;�9- ���1J�.��:]���{���Ѫm5T�M�2`�S���]����Շ����f�"|c�����O���BMG�D���X��s�S�N���=�NH���~�ħC���J.v�i2}	�S�rR��)����8���ر�EGK8��4�ϛ7�(��ͤg�;�z��Y�u���:Y<ͫ'Z�3�Ż�v�*H��b��nY�E�����͍���Q��̏�7.���#�:Q�z7��IЛ9)Ni5���2?Wq�������)&�RY>��aq�������K����vQ_gY�'4rO���qO+rۣ��93u�zq��U%�i?gOj�4=�;:���&nÞ�f�'i=���$���3yԞ5)L�kЖ9��V�
H�1��Y&��J�6]T�9�=�7��(�w�t�����jn0�Yb���h�g!����ѢǍ*KS%޶�h]F�ɩ�2X��}�b+���'��1'�T��g:p�7��t�C�p{����w��:b���q]e:�؝�͊}gR��Qa��#Eɬ�动;��Ns��?c�<m��9��FE/�t�RR�+S��nغ�Yv�[�nmdM����&e�-M�zZ�3��8&�e2Z�%�v0x�5f�)'��w���q8�y��Hp�)��T�I���/>�LjڲGdɽ��Ne�ɩ���Xxdʔ�)����S��z�I<�*H��M�]��BBl�"�