BZh91AY&SY��o _�Py���������`�       � �`�2��� �`�2��� �`�2��� �`�2��� �`�2��*HAD� M=@z����SM�݀��	`�B4�����b�����F��H��ʓ�^����3T�����RI���y;��*�7�Ś.�*�♼l,�o���rY�w����M�^�����j�L�))z�Y�L3R�v��)��+³nۙ�έlp7.�u���zM4���*��M8�vW����Y�SFצH���a���Hp���M�����c���4�R�UUv�U�#�O�����BΊ�\b�X�nK^��][뢚=S��d��n��kY��H���z����´��U�b燃)���{gm�2�oM^
�߳\��l庰��]cJؼ㥡�%�f/k�S�+6Se-Rl����a���c�R͆Q},�K���y+]�/j^�o�-�e����G��i���ʪ�YQ�x�����r�JR�\UUUUUT�*ʞ�����<`��G�M�y�R�Qg�=+���,�Ҳ�����V0��3�-�eP�kJŭUl^��ҔMer���mT�SmO[j�-E��zvR�)F�M�W�/u���g��ϖ�_;��8S��d�\Z�/w�vʹ���X�K���S��O��Si��2lY�j��U��Z텎�f�=N����{�>���<�����a��̍G�C�AcЍ�"���n~����a�,��9�.��Qs�H��O�8�~Ε)L"�:�#��'�[�Z���R�>L���Ee�m#<�{��U��7.�x{�C'�ڲxa��--�v.d�"��Ja�fm.��;����QgqG��A���H��d�<�Q�y�7��$�M�*S����r�����a�}��~\�#GL�O9y0�(�d�#��OZbS�vrX���#���0�p���16=�I�n[tvgK7P��IʑeRX���r�m_��F��G_�?��f�9����w���(�x��U'r���i�y��38j�aIC�8,�%rR�Y�JS��ڱ�z�M�Qt���/��)�40ݰ�
ae�*G�Z<�3&��h�c�*KS%ަ�h]F�ɩ��cW������C�{�eI)�9���ܺO�������6�gD]#���K��;�:ӝw[��O9ԩ#�Xw����q��㊨:���9���9��h�7�������UE/�l�RR�+S��d]GK.σsb�ͬ��#���Jf]x�6m�j38���of�2Z�s���%�u�xx�f�]MT�8����`g�G���T���
�H��/<��յd�C&M��tt�1;��&T�rLgF�ƝE;�ZI�QRF��h���H�
�-�