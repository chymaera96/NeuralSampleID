BZh91AY&SY3�� _�Py���������`� @    `�1 �&	�!��L��`�1 �&	�!��L���{M4  h  � �0L@0	�h�h`bc�0L@0	�h�h`b`�"2�=h�i�G���i7aw�KHLa��g괆R���(�Q*�D�*O�z���K�2T��R2P1��:O��W����E��
dɂ���E��+;.��9�T�l�`��)*y�kL��1S;������޳��2��cyuۗ]���'�Yy��J�<^�,�L��\ŷFk�z����3a��#D�&��G��W�Y&��
�����v��Q��P����_َ*����u��v�W����5eL}s�b�f��Wi)��URl��U��UUD*���ng���7R��=Y6�>T��i17,���7�6�*�e:�u������CP��	�3Hl	(�Ą�)ajjd2��̳�X�͗eg8Suߖ5�k�߫L�ڳ��V\��7��ն�lnZ]������x*��)U�UUUUUUIP������;�|T�OAJQe~�H�.�f,��-f�j��Vv�U�j�&Y�0M�fɑ�cj�n��&ʑJmF3��vlV�����G5�u&�/w�\>�_L�v����������],_ϡ���>+�ښ9;�	v�w�}O���D��R��Y��N���>�]�c������=�7���ǝ=i>6d>i*��E���F�Obu7?$���9���,��N�7��(��$|���'O��JSSg]$rE���"ڨu2���K,���
H���&q�P�q:*�Qf��/�:��V�'c�cp�i�Tb�"�$
J`ܳ6k`��̅�["���䘟n-j����s�J:����>�'Jk�Jp�I��Q���;�������*FnrY=��q�����N}���"줱7]�G'�����9������'�ܶ��<���:�ɽ9T�*�ų�����e�Y�f{�v�Gങ;N��������'�IG[�2yԞ
R:�&ϙ,t2��L���)�i%rR�Y���Eǹc�I&�(�x�u������47)��,Q?����C)F�5��-L%޶ih]F�š�1X��|�"+��퇵�0���IO�МH޾��|O�������}k:����r]e:]	ڝ+�]�T�j�=E���܌׆�'�Pv�ö���П7c{c���p�8#QKĩ�;Ԕ�����gc�.��=�{sU�1&���Ly�E�-Mv�i�.���1Rʳ��Ĥ�����FN����y�W}m0D���d��!��R�T��<���`uF��H�X��g#�����w;��,iH�eFg��e<VZI�QRF�����ܑN$� � 