BZh91AY&SYϡ�� ;߀Py���������`�T���   9�#� �&���0F&9�#� �&���0F&9�#� �&���0F&�"jh����h42  hM 9�#� �&���0F&
� �b24�@L
P6�'��57�5�!]QГ���������d��0TJ�RH��,�>��W�$���R#�H�H1��:N���ګ~n��\n�Č$q����It�6���X�D�	�SH�dn��IEgr
��	��س>{�L�}6��6.�d䪱�h��	`��r0X���NϾ`0k��T�l�V�/�CdiN�й�����ʬS9�UU����8��Q��)����0oȇf�)Sz�F�QTD��Z�w��(��"sfa ��w���
����3��ʓU"��L�e)�Kƚ���ا���P�PEGh�-�VڳrI0n`����i%h��b��K��[Ŋ��=,ʄK!����#��j�O��������ɪ���J&U�#%w|
�w����)j\�3Q$�!9#�h7!��!-�$�J����Yi����4`Yң�R5Jy�q�@����$dI28��:n���3$��;�L�@$ ��\��,Ft�Y�I�R)MTc=M+�b��!�<�l@�2f��" �<���eɺ���T��X������]�U47�K��Fwa3ݰ�q���C�$6��Is�<9�40y�^��#i>Q����O/Ğ�X�j�}"�X�[ȧ�9��D��"�a��r)���}�.t���	�S��)�)����7���VqV̣�祖~���
H���&q�R;�M�X��Z�����^6���6)u�N���ҲE�pb))�Z̙�]���24�"���1<$k-j�����(�<�D�I9SO)�M'�F"���`�=��~;\��D��K'���#�w1{��NS	M��Ibk���WA��dpN�	��oOZ���4�d瑽ț�%�Ib��ݼS��~Vlٞ�z#�ZL�M� �N�9�Q��;ԝ�R9�&��,ne&
H�a�شL��J�4�T�7\z�1���(�wh9���|�d��f
`����Z:He#Ta�X�J����]�f���hV-r1X��{"+���G���I�$���6�r/�t����kI��,拤q;���S��8�*�.��<�:��Aa��kFk��"x��/X�#q�������3t9�K\pc،E/�T�RR�+A�r·L]Gz~Mm*5�1&�N�&<"떦�\�26�&��1Z��V�Ғ�8�:��2r�����w��s�M�ݬ��Hm�Sc�R*'�Iy�09�CR��b����&�����t��\Xґ�0ʌϝ9�w,���EI\����ܑN$3�v~�